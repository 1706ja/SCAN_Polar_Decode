module opcode #(parameter P = 32) (clk, rst, channel, I_program_counter,O_opcode, O_opcode_next, O_opcode_delay,
        O_Nv,O_Nv_next, O_part_count,O_part_count_next, O_address, O_address_next, O_opcode_before, O_Nv_before, O_bit_count);
        input clk,rst;
        input channel;
        input [15:0] I_program_counter;
        output [3:0] O_opcode,O_opcode_next, O_opcode_before, O_opcode_delay;
        output [10:0] O_Nv, O_Nv_next, O_Nv_before;
        output [4:0] O_part_count, O_part_count_next;
        output [9:0] O_address, O_address_next;
        output [12:0] O_bit_count;
        localparam TYPE1     = 4'b0000;
        localparam TYPE2     = 4'b0001;
        localparam BOTTOM    = 4'b0010;
        localparam TYPE3     = 4'b0011;
        localparam IDLE      = 4'b1011;

        reg [3:0] L_opcode, L_opcode_next, L_opcode_before, L_opcode_delay;
        reg [10:0] L_Nv,L_Nv_next,L_Nv_before, L_Nv_delay;
        reg [4:0] L_part_count, L_part_count_next, L_part_count_delay;
        reg [9:0] Address, Address_next, Address_delay;
        reg[12:0] L_bit_count;
        
        // assignment of outputs
        assign O_opcode = L_opcode;
        assign O_opcode_delay = L_opcode_delay;
        assign O_opcode_next = L_opcode_next;
        assign O_opcode_before = L_opcode_before;
        assign O_Nv = L_Nv;
        assign O_Nv_next = L_Nv_next;
        assign O_Nv_before = L_Nv_before;
        assign O_part_count = L_part_count;
        assign O_part_count_next = L_part_count_next;
        assign O_address = Address;
        assign O_address_next = Address_next;
        assign O_bit_count = L_bit_count;


        wire islast, oprand;
       assign islast = (L_Nv_next) > (2*P*(1+L_part_count_next));
       assign oprand = (L_opcode_next==TYPE1||L_opcode_next==TYPE2);

       always @(posedge clk)
     begin       
           if(!rst) begin
                L_Nv_before <= L_Nv;        
                L_Nv <= L_Nv_delay;
                L_Nv_delay <= L_Nv_next;

                L_opcode_before <= L_opcode;
                L_opcode <= L_opcode_delay;
                L_opcode_delay <= L_opcode_next;


                L_part_count <= L_part_count_delay;
                L_part_count_delay <= L_part_count_next;

//                Address_before <= Address;       
                L_bit_count <= (L_bit_count+2*(L_opcode==BOTTOM));

                Address <= Address_delay;
                Address_delay <= Address_next;
            end
            else begin
              L_bit_count <= 0;
              L_Nv                          <=1024; 
              L_Nv_before                          <=1024; 
              L_Nv_delay                          <=1024; 

              L_opcode_before <= TYPE1;
              L_opcode <= TYPE1;
              L_opcode_delay <= TYPE1;


              L_part_count <= 0;
              L_part_count_delay <= 0;

              Address <= 0;
              Address_delay <= 0;
            end
        end



        always @(posedge clk) begin
            if(rst) begin
            
            L_Nv_next                     <=1024;
            L_opcode_next <= TYPE1;
            L_part_count_next <= 0;
            // Address <= -1;
            Address_next <= 0;
            end
            else begin
           if (channel) begin
              case (L_Nv_next)
                1024 : L_Nv_next <= islast ? 1024 : 512;
                512 : L_Nv_next <= islast ?  512 : (oprand?256:1024);
                256 : L_Nv_next <= islast ? 256 : (oprand?128:512);
                128 : L_Nv_next <= oprand ? 64 : 256;
                64 : L_Nv_next <= oprand ? 32 : 128;
                32 : L_Nv_next <= oprand ? 16 : 64;
                16 : L_Nv_next <= oprand ? 8 : 32;
                8 : L_Nv_next <= oprand ? 4 : 16;
                4 : L_Nv_next <= oprand ? 2 : 8;
                2 : L_Nv_next <= 4;
                default: L_Nv_next <= 1024;
              endcase

              case (L_opcode_next)
                TYPE1 : L_opcode_next <= islast ? TYPE1 : ( (L_Nv_next==4) ? BOTTOM : TYPE1 );
                TYPE2 : L_opcode_next <= islast ? TYPE2 : ( (L_Nv_next==4) ? BOTTOM : TYPE1 );
                TYPE3 : L_opcode_next <= islast ? TYPE3 : ( (Address_next[0]) ? TYPE3 : TYPE2);
                BOTTOM : L_opcode_next <= Address_next[0] ? TYPE3 : TYPE2 ;
                default: L_opcode_next <= TYPE1;
              endcase

                // case (L_part_count_next)
                //   0 : L_part_count_next <= (L_Nv_next>2*P) ? 1 : 0;
                //   1 : L_part_count_next <= (L_Nv_next>4*P) ? 2 : 0;
                //   2 : L_part_count_next <= (L_Nv_next>4*P) ? 3 : 0;
                //   3 : L_part_count_next <=  0;
                //   4 : L_part_count_next <= (L_Nv_next>8*P) ? 5 : 0;
                //   5 : L_part_count_next <= (L_Nv_next>8*P) ? 6 : 0;
                //   6 : L_part_count_next <= (L_Nv_next>8*P) ? 7 : 0;
                //   7 : L_part_count_next <= 0;
                //   default: L_part_count_next <= 0;
                // endcase
                L_part_count_next <= islast ? (L_part_count_next+1) : 0;


          


      case(I_program_counter)
          34 : Address_next<= 1 ;
          37 : Address_next<= 1 ;
          38 : Address_next<= 2 ;
          40 : Address_next<= 3 ;
          41 : Address_next<= 1 ;
          44 : Address_next<= 1 ;
          45 : Address_next<= 2 ;
          46 : Address_next<= 4 ;
          48 : Address_next<= 5 ;
          49 : Address_next<= 2 ;
          51 : Address_next<= 3 ;
          52 : Address_next<= 6 ;
          54 : Address_next<= 7 ;
          55 : Address_next<= 3 ;
          56 : Address_next<= 1 ;
          59 : Address_next<= 1 ;
          60 : Address_next<= 2 ;
          61 : Address_next<= 4 ;
          62 : Address_next<= 8 ;
          64 : Address_next<= 9 ;
          65 : Address_next<= 4 ;
          67 : Address_next<= 5 ;
          68 : Address_next<= 10 ;
          70 : Address_next<= 11 ;
          71 : Address_next<= 5 ;
          72 : Address_next<= 2 ;
          74 : Address_next<= 3 ;
          75 : Address_next<= 6 ;
          76 : Address_next<= 12 ;
          78 : Address_next<= 13 ;
          79 : Address_next<= 6 ;
          81 : Address_next<= 7 ;
          82 : Address_next<= 14 ;
          84 : Address_next<= 15 ;
          85 : Address_next<= 7 ;
          86 : Address_next<= 3 ;
          87 : Address_next<= 1 ;
          90 : Address_next<= 1 ;
          91 : Address_next<= 2 ;
          92 : Address_next<= 4 ;
          93 : Address_next<= 8 ;
          94 : Address_next<= 16 ;
          96 : Address_next<= 17 ;
          97 : Address_next<= 8 ;
          99 : Address_next<= 9 ;
          100 : Address_next<= 18 ;
          102 : Address_next<= 19 ;
          103 : Address_next<= 9 ;
          104 : Address_next<= 4 ;
          106 : Address_next<= 5 ;
          107 : Address_next<= 10 ;
          108 : Address_next<= 20 ;
          110 : Address_next<= 21 ;
          111 : Address_next<= 10 ;
          113 : Address_next<= 11 ;
          114 : Address_next<= 22 ;
          116 : Address_next<= 23 ;
          117 : Address_next<= 11 ;
          118 : Address_next<= 5 ;
          119 : Address_next<= 2 ;
          121 : Address_next<= 3 ;
          122 : Address_next<= 6 ;
          123 : Address_next<= 12 ;
          124 : Address_next<= 24 ;
          126 : Address_next<= 25 ;
          127 : Address_next<= 12 ;
          129 : Address_next<= 13 ;
          130 : Address_next<= 26 ;
          132 : Address_next<= 27 ;
          133 : Address_next<= 13 ;
          134 : Address_next<= 6 ;
          136 : Address_next<= 7 ;
          137 : Address_next<= 14 ;
          138 : Address_next<= 28 ;
          140 : Address_next<= 29 ;
          141 : Address_next<= 14 ;
          143 : Address_next<= 15 ;
          144 : Address_next<= 30 ;
          146 : Address_next<= 31 ;
          147 : Address_next<= 15 ;
          148 : Address_next<= 7 ;
          149 : Address_next<= 3 ;
          150 : Address_next<= 1 ;
          154 : Address_next<= 1 ;
          155 : Address_next<= 2 ;
          156 : Address_next<= 4 ;
          157 : Address_next<= 8 ;
          158 : Address_next<= 16 ;
          159 : Address_next<= 32 ;
          161 : Address_next<= 33 ;
          162 : Address_next<= 16 ;
          164 : Address_next<= 17 ;
          165 : Address_next<= 34 ;
          167 : Address_next<= 35 ;
          168 : Address_next<= 17 ;
          169 : Address_next<= 8 ;
          171 : Address_next<= 9 ;
          172 : Address_next<= 18 ;
          173 : Address_next<= 36 ;
          175 : Address_next<= 37 ;
          176 : Address_next<= 18 ;
          178 : Address_next<= 19 ;
          179 : Address_next<= 38 ;
          181 : Address_next<= 39 ;
          182 : Address_next<= 19 ;
          183 : Address_next<= 9 ;
          184 : Address_next<= 4 ;
          186 : Address_next<= 5 ;
          187 : Address_next<= 10 ;
          188 : Address_next<= 20 ;
          189 : Address_next<= 40 ;
          191 : Address_next<= 41 ;
          192 : Address_next<= 20 ;
          194 : Address_next<= 21 ;
          195 : Address_next<= 42 ;
          197 : Address_next<= 43 ;
          198 : Address_next<= 21 ;
          199 : Address_next<= 10 ;
          201 : Address_next<= 11 ;
          202 : Address_next<= 22 ;
          203 : Address_next<= 44 ;
          205 : Address_next<= 45 ;
          206 : Address_next<= 22 ;
          208 : Address_next<= 23 ;
          209 : Address_next<= 46 ;
          211 : Address_next<= 47 ;
          212 : Address_next<= 23 ;
          213 : Address_next<= 11 ;
          214 : Address_next<= 5 ;
          215 : Address_next<= 2 ;
          217 : Address_next<= 3 ;
          218 : Address_next<= 6 ;
          219 : Address_next<= 12 ;
          220 : Address_next<= 24 ;
          221 : Address_next<= 48 ;
          223 : Address_next<= 49 ;
          224 : Address_next<= 24 ;
          226 : Address_next<= 25 ;
          227 : Address_next<= 50 ;
          229 : Address_next<= 51 ;
          230 : Address_next<= 25 ;
          231 : Address_next<= 12 ;
          233 : Address_next<= 13 ;
          234 : Address_next<= 26 ;
          235 : Address_next<= 52 ;
          237 : Address_next<= 53 ;
          238 : Address_next<= 26 ;
          240 : Address_next<= 27 ;
          241 : Address_next<= 54 ;
          243 : Address_next<= 55 ;
          244 : Address_next<= 27 ;
          245 : Address_next<= 13 ;
          246 : Address_next<= 6 ;
          248 : Address_next<= 7 ;
          249 : Address_next<= 14 ;
          250 : Address_next<= 28 ;
          251 : Address_next<= 56 ;
          253 : Address_next<= 57 ;
          254 : Address_next<= 28 ;
          256 : Address_next<= 29 ;
          257 : Address_next<= 58 ;
          259 : Address_next<= 59 ;
          260 : Address_next<= 29 ;
          261 : Address_next<= 14 ;
          263 : Address_next<= 15 ;
          264 : Address_next<= 30 ;
          265 : Address_next<= 60 ;
          267 : Address_next<= 61 ;
          268 : Address_next<= 30 ;
          270 : Address_next<= 31 ;
          271 : Address_next<= 62 ;
          273 : Address_next<= 63 ;
          274 : Address_next<= 31 ;
          275 : Address_next<= 15 ;
          276 : Address_next<= 7 ;
          277 : Address_next<= 3 ;
          278 : Address_next<= 1 ;
          285 : Address_next<= 1 ;
          286 : Address_next<= 1 ;
          287 : Address_next<= 2 ;
          288 : Address_next<= 4 ;
          289 : Address_next<= 8 ;
          290 : Address_next<= 16 ;
          291 : Address_next<= 32 ;
          292 : Address_next<= 64 ;
          294 : Address_next<= 65 ;
          295 : Address_next<= 32 ;
          297 : Address_next<= 33 ;
          298 : Address_next<= 66 ;
          300 : Address_next<= 67 ;
          301 : Address_next<= 33 ;
          302 : Address_next<= 16 ;
          304 : Address_next<= 17 ;
          305 : Address_next<= 34 ;
          306 : Address_next<= 68 ;
          308 : Address_next<= 69 ;
          309 : Address_next<= 34 ;
          311 : Address_next<= 35 ;
          312 : Address_next<= 70 ;
          314 : Address_next<= 71 ;
          315 : Address_next<= 35 ;
          316 : Address_next<= 17 ;
          317 : Address_next<= 8 ;
          319 : Address_next<= 9 ;
          320 : Address_next<= 18 ;
          321 : Address_next<= 36 ;
          322 : Address_next<= 72 ;
          324 : Address_next<= 73 ;
          325 : Address_next<= 36 ;
          327 : Address_next<= 37 ;
          328 : Address_next<= 74 ;
          330 : Address_next<= 75 ;
          331 : Address_next<= 37 ;
          332 : Address_next<= 18 ;
          334 : Address_next<= 19 ;
          335 : Address_next<= 38 ;
          336 : Address_next<= 76 ;
          338 : Address_next<= 77 ;
          339 : Address_next<= 38 ;
          341 : Address_next<= 39 ;
          342 : Address_next<= 78 ;
          344 : Address_next<= 79 ;
          345 : Address_next<= 39 ;
          346 : Address_next<= 19 ;
          347 : Address_next<= 9 ;
          348 : Address_next<= 4 ;
          350 : Address_next<= 5 ;
          351 : Address_next<= 10 ;
          352 : Address_next<= 20 ;
          353 : Address_next<= 40 ;
          354 : Address_next<= 80 ;
          356 : Address_next<= 81 ;
          357 : Address_next<= 40 ;
          359 : Address_next<= 41 ;
          360 : Address_next<= 82 ;
          362 : Address_next<= 83 ;
          363 : Address_next<= 41 ;
          364 : Address_next<= 20 ;
          366 : Address_next<= 21 ;
          367 : Address_next<= 42 ;
          368 : Address_next<= 84 ;
          370 : Address_next<= 85 ;
          371 : Address_next<= 42 ;
          373 : Address_next<= 43 ;
          374 : Address_next<= 86 ;
          376 : Address_next<= 87 ;
          377 : Address_next<= 43 ;
          378 : Address_next<= 21 ;
          379 : Address_next<= 10 ;
          381 : Address_next<= 11 ;
          382 : Address_next<= 22 ;
          383 : Address_next<= 44 ;
          384 : Address_next<= 88 ;
          386 : Address_next<= 89 ;
          387 : Address_next<= 44 ;
          389 : Address_next<= 45 ;
          390 : Address_next<= 90 ;
          392 : Address_next<= 91 ;
          393 : Address_next<= 45 ;
          394 : Address_next<= 22 ;
          396 : Address_next<= 23 ;
          397 : Address_next<= 46 ;
          398 : Address_next<= 92 ;
          400 : Address_next<= 93 ;
          401 : Address_next<= 46 ;
          403 : Address_next<= 47 ;
          404 : Address_next<= 94 ;
          406 : Address_next<= 95 ;
          407 : Address_next<= 47 ;
          408 : Address_next<= 23 ;
          409 : Address_next<= 11 ;
          410 : Address_next<= 5 ;
          411 : Address_next<= 2 ;
          414 : Address_next<= 3 ;
          415 : Address_next<= 6 ;
          416 : Address_next<= 12 ;
          417 : Address_next<= 24 ;
          418 : Address_next<= 48 ;
          419 : Address_next<= 96 ;
          421 : Address_next<= 97 ;
          422 : Address_next<= 48 ;
          424 : Address_next<= 49 ;
          425 : Address_next<= 98 ;
          427 : Address_next<= 99 ;
          428 : Address_next<= 49 ;
          429 : Address_next<= 24 ;
          431 : Address_next<= 25 ;
          432 : Address_next<= 50 ;
          433 : Address_next<= 100 ;
          435 : Address_next<= 101 ;
          436 : Address_next<= 50 ;
          438 : Address_next<= 51 ;
          439 : Address_next<= 102 ;
          441 : Address_next<= 103 ;
          442 : Address_next<= 51 ;
          443 : Address_next<= 25 ;
          444 : Address_next<= 12 ;
          446 : Address_next<= 13 ;
          447 : Address_next<= 26 ;
          448 : Address_next<= 52 ;
          449 : Address_next<= 104 ;
          451 : Address_next<= 105 ;
          452 : Address_next<= 52 ;
          454 : Address_next<= 53 ;
          455 : Address_next<= 106 ;
          457 : Address_next<= 107 ;
          458 : Address_next<= 53 ;
          459 : Address_next<= 26 ;
          461 : Address_next<= 27 ;
          462 : Address_next<= 54 ;
          463 : Address_next<= 108 ;
          465 : Address_next<= 109 ;
          466 : Address_next<= 54 ;
          468 : Address_next<= 55 ;
          469 : Address_next<= 110 ;
          471 : Address_next<= 111 ;
          472 : Address_next<= 55 ;
          473 : Address_next<= 27 ;
          474 : Address_next<= 13 ;
          475 : Address_next<= 6 ;
          477 : Address_next<= 7 ;
          478 : Address_next<= 14 ;
          479 : Address_next<= 28 ;
          480 : Address_next<= 56 ;
          481 : Address_next<= 112 ;
          483 : Address_next<= 113 ;
          484 : Address_next<= 56 ;
          486 : Address_next<= 57 ;
          487 : Address_next<= 114 ;
          489 : Address_next<= 115 ;
          490 : Address_next<= 57 ;
          491 : Address_next<= 28 ;
          493 : Address_next<= 29 ;
          494 : Address_next<= 58 ;
          495 : Address_next<= 116 ;
          497 : Address_next<= 117 ;
          498 : Address_next<= 58 ;
          500 : Address_next<= 59 ;
          501 : Address_next<= 118 ;
          503 : Address_next<= 119 ;
          504 : Address_next<= 59 ;
          505 : Address_next<= 29 ;
          506 : Address_next<= 14 ;
          508 : Address_next<= 15 ;
          509 : Address_next<= 30 ;
          510 : Address_next<= 60 ;
          511 : Address_next<= 120 ;
          513 : Address_next<= 121 ;
          514 : Address_next<= 60 ;
          516 : Address_next<= 61 ;
          517 : Address_next<= 122 ;
          519 : Address_next<= 123 ;
          520 : Address_next<= 61 ;
          521 : Address_next<= 30 ;
          523 : Address_next<= 31 ;
          524 : Address_next<= 62 ;
          525 : Address_next<= 124 ;
          527 : Address_next<= 125 ;
          528 : Address_next<= 62 ;
          530 : Address_next<= 63 ;
          531 : Address_next<= 126 ;
          533 : Address_next<= 127 ;
          534 : Address_next<= 63 ;
          535 : Address_next<= 31 ;
          536 : Address_next<= 15 ;
          537 : Address_next<= 7 ;
          538 : Address_next<= 3 ;
          539 : Address_next<= 1 ;
          540 : Address_next<= 1 ;
          553 : Address_next<= 1 ;
          554 : Address_next<= 1 ;
          555 : Address_next<= 1 ;
          556 : Address_next<= 1 ;
          557 : Address_next<= 2 ;
          558 : Address_next<= 2 ;
          559 : Address_next<= 4 ;
          560 : Address_next<= 8 ;
          561 : Address_next<= 16 ;
          562 : Address_next<= 32 ;
          563 : Address_next<= 64 ;
          564 : Address_next<= 128 ;
          566 : Address_next<= 129 ;
          567 : Address_next<= 64 ;
          569 : Address_next<= 65 ;
          570 : Address_next<= 130 ;
          572 : Address_next<= 131 ;
          573 : Address_next<= 65 ;
          574 : Address_next<= 32 ;
          576 : Address_next<= 33 ;
          577 : Address_next<= 66 ;
          578 : Address_next<= 132 ;
          580 : Address_next<= 133 ;
          581 : Address_next<= 66 ;
          583 : Address_next<= 67 ;
          584 : Address_next<= 134 ;
          586 : Address_next<= 135 ;
          587 : Address_next<= 67 ;
          588 : Address_next<= 33 ;
          589 : Address_next<= 16 ;
          591 : Address_next<= 17 ;
          592 : Address_next<= 34 ;
          593 : Address_next<= 68 ;
          594 : Address_next<= 136 ;
          596 : Address_next<= 137 ;
          597 : Address_next<= 68 ;
          599 : Address_next<= 69 ;
          600 : Address_next<= 138 ;
          602 : Address_next<= 139 ;
          603 : Address_next<= 69 ;
          604 : Address_next<= 34 ;
          606 : Address_next<= 35 ;
          607 : Address_next<= 70 ;
          608 : Address_next<= 140 ;
          610 : Address_next<= 141 ;
          611 : Address_next<= 70 ;
          613 : Address_next<= 71 ;
          614 : Address_next<= 142 ;
          616 : Address_next<= 143 ;
          617 : Address_next<= 71 ;
          618 : Address_next<= 35 ;
          619 : Address_next<= 17 ;
          620 : Address_next<= 8 ;
          622 : Address_next<= 9 ;
          623 : Address_next<= 18 ;
          624 : Address_next<= 36 ;
          625 : Address_next<= 72 ;
          626 : Address_next<= 144 ;
          628 : Address_next<= 145 ;
          629 : Address_next<= 72 ;
          631 : Address_next<= 73 ;
          632 : Address_next<= 146 ;
          634 : Address_next<= 147 ;
          635 : Address_next<= 73 ;
          636 : Address_next<= 36 ;
          638 : Address_next<= 37 ;
          639 : Address_next<= 74 ;
          640 : Address_next<= 148 ;
          642 : Address_next<= 149 ;
          643 : Address_next<= 74 ;
          645 : Address_next<= 75 ;
          646 : Address_next<= 150 ;
          648 : Address_next<= 151 ;
          649 : Address_next<= 75 ;
          650 : Address_next<= 37 ;
          651 : Address_next<= 18 ;
          653 : Address_next<= 19 ;
          654 : Address_next<= 38 ;
          655 : Address_next<= 76 ;
          656 : Address_next<= 152 ;
          658 : Address_next<= 153 ;
          659 : Address_next<= 76 ;
          661 : Address_next<= 77 ;
          662 : Address_next<= 154 ;
          664 : Address_next<= 155 ;
          665 : Address_next<= 77 ;
          666 : Address_next<= 38 ;
          668 : Address_next<= 39 ;
          669 : Address_next<= 78 ;
          670 : Address_next<= 156 ;
          672 : Address_next<= 157 ;
          673 : Address_next<= 78 ;
          675 : Address_next<= 79 ;
          676 : Address_next<= 158 ;
          678 : Address_next<= 159 ;
          679 : Address_next<= 79 ;
          680 : Address_next<= 39 ;
          681 : Address_next<= 19 ;
          682 : Address_next<= 9 ;
          683 : Address_next<= 4 ;
          686 : Address_next<= 5 ;
          687 : Address_next<= 10 ;
          688 : Address_next<= 20 ;
          689 : Address_next<= 40 ;
          690 : Address_next<= 80 ;
          691 : Address_next<= 160 ;
          693 : Address_next<= 161 ;
          694 : Address_next<= 80 ;
          696 : Address_next<= 81 ;
          697 : Address_next<= 162 ;
          699 : Address_next<= 163 ;
          700 : Address_next<= 81 ;
          701 : Address_next<= 40 ;
          703 : Address_next<= 41 ;
          704 : Address_next<= 82 ;
          705 : Address_next<= 164 ;
          707 : Address_next<= 165 ;
          708 : Address_next<= 82 ;
          710 : Address_next<= 83 ;
          711 : Address_next<= 166 ;
          713 : Address_next<= 167 ;
          714 : Address_next<= 83 ;
          715 : Address_next<= 41 ;
          716 : Address_next<= 20 ;
          718 : Address_next<= 21 ;
          719 : Address_next<= 42 ;
          720 : Address_next<= 84 ;
          721 : Address_next<= 168 ;
          723 : Address_next<= 169 ;
          724 : Address_next<= 84 ;
          726 : Address_next<= 85 ;
          727 : Address_next<= 170 ;
          729 : Address_next<= 171 ;
          730 : Address_next<= 85 ;
          731 : Address_next<= 42 ;
          733 : Address_next<= 43 ;
          734 : Address_next<= 86 ;
          735 : Address_next<= 172 ;
          737 : Address_next<= 173 ;
          738 : Address_next<= 86 ;
          740 : Address_next<= 87 ;
          741 : Address_next<= 174 ;
          743 : Address_next<= 175 ;
          744 : Address_next<= 87 ;
          745 : Address_next<= 43 ;
          746 : Address_next<= 21 ;
          747 : Address_next<= 10 ;
          749 : Address_next<= 11 ;
          750 : Address_next<= 22 ;
          751 : Address_next<= 44 ;
          752 : Address_next<= 88 ;
          753 : Address_next<= 176 ;
          755 : Address_next<= 177 ;
          756 : Address_next<= 88 ;
          758 : Address_next<= 89 ;
          759 : Address_next<= 178 ;
          761 : Address_next<= 179 ;
          762 : Address_next<= 89 ;
          763 : Address_next<= 44 ;
          765 : Address_next<= 45 ;
          766 : Address_next<= 90 ;
          767 : Address_next<= 180 ;
          769 : Address_next<= 181 ;
          770 : Address_next<= 90 ;
          772 : Address_next<= 91 ;
          773 : Address_next<= 182 ;
          775 : Address_next<= 183 ;
          776 : Address_next<= 91 ;
          777 : Address_next<= 45 ;
          778 : Address_next<= 22 ;
          780 : Address_next<= 23 ;
          781 : Address_next<= 46 ;
          782 : Address_next<= 92 ;
          783 : Address_next<= 184 ;
          785 : Address_next<= 185 ;
          786 : Address_next<= 92 ;
          788 : Address_next<= 93 ;
          789 : Address_next<= 186 ;
          791 : Address_next<= 187 ;
          792 : Address_next<= 93 ;
          793 : Address_next<= 46 ;
          795 : Address_next<= 47 ;
          796 : Address_next<= 94 ;
          797 : Address_next<= 188 ;
          799 : Address_next<= 189 ;
          800 : Address_next<= 94 ;
          802 : Address_next<= 95 ;
          803 : Address_next<= 190 ;
          805 : Address_next<= 191 ;
          806 : Address_next<= 95 ;
          807 : Address_next<= 47 ;
          808 : Address_next<= 23 ;
          809 : Address_next<= 11 ;
          810 : Address_next<= 5 ;
          811 : Address_next<= 2 ;
          812 : Address_next<= 2 ;
          817 : Address_next<= 3 ;
          818 : Address_next<= 3 ;
          819 : Address_next<= 6 ;
          820 : Address_next<= 12 ;
          821 : Address_next<= 24 ;
          822 : Address_next<= 48 ;
          823 : Address_next<= 96 ;
          824 : Address_next<= 192 ;
          826 : Address_next<= 193 ;
          827 : Address_next<= 96 ;
          829 : Address_next<= 97 ;
          830 : Address_next<= 194 ;
          832 : Address_next<= 195 ;
          833 : Address_next<= 97 ;
          834 : Address_next<= 48 ;
          836 : Address_next<= 49 ;
          837 : Address_next<= 98 ;
          838 : Address_next<= 196 ;
          840 : Address_next<= 197 ;
          841 : Address_next<= 98 ;
          843 : Address_next<= 99 ;
          844 : Address_next<= 198 ;
          846 : Address_next<= 199 ;
          847 : Address_next<= 99 ;
          848 : Address_next<= 49 ;
          849 : Address_next<= 24 ;
          851 : Address_next<= 25 ;
          852 : Address_next<= 50 ;
          853 : Address_next<= 100 ;
          854 : Address_next<= 200 ;
          856 : Address_next<= 201 ;
          857 : Address_next<= 100 ;
          859 : Address_next<= 101 ;
          860 : Address_next<= 202 ;
          862 : Address_next<= 203 ;
          863 : Address_next<= 101 ;
          864 : Address_next<= 50 ;
          866 : Address_next<= 51 ;
          867 : Address_next<= 102 ;
          868 : Address_next<= 204 ;
          870 : Address_next<= 205 ;
          871 : Address_next<= 102 ;
          873 : Address_next<= 103 ;
          874 : Address_next<= 206 ;
          876 : Address_next<= 207 ;
          877 : Address_next<= 103 ;
          878 : Address_next<= 51 ;
          879 : Address_next<= 25 ;
          880 : Address_next<= 12 ;
          882 : Address_next<= 13 ;
          883 : Address_next<= 26 ;
          884 : Address_next<= 52 ;
          885 : Address_next<= 104 ;
          886 : Address_next<= 208 ;
          888 : Address_next<= 209 ;
          889 : Address_next<= 104 ;
          891 : Address_next<= 105 ;
          892 : Address_next<= 210 ;
          894 : Address_next<= 211 ;
          895 : Address_next<= 105 ;
          896 : Address_next<= 52 ;
          898 : Address_next<= 53 ;
          899 : Address_next<= 106 ;
          900 : Address_next<= 212 ;
          902 : Address_next<= 213 ;
          903 : Address_next<= 106 ;
          905 : Address_next<= 107 ;
          906 : Address_next<= 214 ;
          908 : Address_next<= 215 ;
          909 : Address_next<= 107 ;
          910 : Address_next<= 53 ;
          911 : Address_next<= 26 ;
          913 : Address_next<= 27 ;
          914 : Address_next<= 54 ;
          915 : Address_next<= 108 ;
          916 : Address_next<= 216 ;
          918 : Address_next<= 217 ;
          919 : Address_next<= 108 ;
          921 : Address_next<= 109 ;
          922 : Address_next<= 218 ;
          924 : Address_next<= 219 ;
          925 : Address_next<= 109 ;
          926 : Address_next<= 54 ;
          928 : Address_next<= 55 ;
          929 : Address_next<= 110 ;
          930 : Address_next<= 220 ;
          932 : Address_next<= 221 ;
          933 : Address_next<= 110 ;
          935 : Address_next<= 111 ;
          936 : Address_next<= 222 ;
          938 : Address_next<= 223 ;
          939 : Address_next<= 111 ;
          940 : Address_next<= 55 ;
          941 : Address_next<= 27 ;
          942 : Address_next<= 13 ;
          943 : Address_next<= 6 ;
          946 : Address_next<= 7 ;
          947 : Address_next<= 14 ;
          948 : Address_next<= 28 ;
          949 : Address_next<= 56 ;
          950 : Address_next<= 112 ;
          951 : Address_next<= 224 ;
          953 : Address_next<= 225 ;
          954 : Address_next<= 112 ;
          956 : Address_next<= 113 ;
          957 : Address_next<= 226 ;
          959 : Address_next<= 227 ;
          960 : Address_next<= 113 ;
          961 : Address_next<= 56 ;
          963 : Address_next<= 57 ;
          964 : Address_next<= 114 ;
          965 : Address_next<= 228 ;
          967 : Address_next<= 229 ;
          968 : Address_next<= 114 ;
          970 : Address_next<= 115 ;
          971 : Address_next<= 230 ;
          973 : Address_next<= 231 ;
          974 : Address_next<= 115 ;
          975 : Address_next<= 57 ;
          976 : Address_next<= 28 ;
          978 : Address_next<= 29 ;
          979 : Address_next<= 58 ;
          980 : Address_next<= 116 ;
          981 : Address_next<= 232 ;
          983 : Address_next<= 233 ;
          984 : Address_next<= 116 ;
          986 : Address_next<= 117 ;
          987 : Address_next<= 234 ;
          989 : Address_next<= 235 ;
          990 : Address_next<= 117 ;
          991 : Address_next<= 58 ;
          993 : Address_next<= 59 ;
          994 : Address_next<= 118 ;
          995 : Address_next<= 236 ;
          997 : Address_next<= 237 ;
          998 : Address_next<= 118 ;
          1000 : Address_next<= 119 ;
          1001 : Address_next<= 238 ;
          1003 : Address_next<= 239 ;
          1004 : Address_next<= 119 ;
          1005 : Address_next<= 59 ;
          1006 : Address_next<= 29 ;
          1007 : Address_next<= 14 ;
          1009 : Address_next<= 15 ;
          1010 : Address_next<= 30 ;
          1011 : Address_next<= 60 ;
          1012 : Address_next<= 120 ;
          1013 : Address_next<= 240 ;
          1015 : Address_next<= 241 ;
          1016 : Address_next<= 120 ;
          1018 : Address_next<= 121 ;
          1019 : Address_next<= 242 ;
          1021 : Address_next<= 243 ;
          1022 : Address_next<= 121 ;
          1023 : Address_next<= 60 ;
          1025 : Address_next<= 61 ;
          1026 : Address_next<= 122 ;
          1027 : Address_next<= 244 ;
          1029 : Address_next<= 245 ;
          1030 : Address_next<= 122 ;
          1032 : Address_next<= 123 ;
          1033 : Address_next<= 246 ;
          1035 : Address_next<= 247 ;
          1036 : Address_next<= 123 ;
          1037 : Address_next<= 61 ;
          1038 : Address_next<= 30 ;
          1040 : Address_next<= 31 ;
          1041 : Address_next<= 62 ;
          1042 : Address_next<= 124 ;
          1043 : Address_next<= 248 ;
          1045 : Address_next<= 249 ;
          1046 : Address_next<= 124 ;
          1048 : Address_next<= 125 ;
          1049 : Address_next<= 250 ;
          1051 : Address_next<= 251 ;
          1052 : Address_next<= 125 ;
          1053 : Address_next<= 62 ;
          1055 : Address_next<= 63 ;
          1056 : Address_next<= 126 ;
          1057 : Address_next<= 252 ;
          1059 : Address_next<= 253 ;
          1060 : Address_next<= 126 ;
          1062 : Address_next<= 127 ;
          1063 : Address_next<= 254 ;
          1065 : Address_next<= 255 ;
          1066 : Address_next<= 127 ;
          1067 : Address_next<= 63 ;
          1068 : Address_next<= 31 ;
          1069 : Address_next<= 15 ;
          1070 : Address_next<= 7 ;
          1071 : Address_next<= 3 ;
          1072 : Address_next<= 3 ;
          1073 : Address_next<= 1 ;
          1074 : Address_next<= 1 ;
          1075 : Address_next<= 1 ;
          1076 : Address_next<= 1 ;
          1101 : Address_next<= 1 ;
          1102 : Address_next<= 1 ;
          1103 : Address_next<= 1 ;
          1104 : Address_next<= 1 ;
          1105 : Address_next<= 1 ;
          1106 : Address_next<= 1 ;
          1107 : Address_next<= 1 ;
          1108 : Address_next<= 1 ;
          1109 : Address_next<= 2 ;
          1110 : Address_next<= 2 ;
          1111 : Address_next<= 2 ;
          1112 : Address_next<= 2 ;
          1113 : Address_next<= 4 ;
          1114 : Address_next<= 4 ;
          1115 : Address_next<= 8 ;
          1116 : Address_next<= 16 ;
          1117 : Address_next<= 32 ;
          1118 : Address_next<= 64 ;
          1119 : Address_next<= 128 ;
          1120 : Address_next<= 256 ;
          1122 : Address_next<= 257 ;
          1123 : Address_next<= 128 ;
          1125 : Address_next<= 129 ;
          1126 : Address_next<= 258 ;
          1128 : Address_next<= 259 ;
          1129 : Address_next<= 129 ;
          1130 : Address_next<= 64 ;
          1132 : Address_next<= 65 ;
          1133 : Address_next<= 130 ;
          1134 : Address_next<= 260 ;
          1136 : Address_next<= 261 ;
          1137 : Address_next<= 130 ;
          1139 : Address_next<= 131 ;
          1140 : Address_next<= 262 ;
          1142 : Address_next<= 263 ;
          1143 : Address_next<= 131 ;
          1144 : Address_next<= 65 ;
          1145 : Address_next<= 32 ;
          1147 : Address_next<= 33 ;
          1148 : Address_next<= 66 ;
          1149 : Address_next<= 132 ;
          1150 : Address_next<= 264 ;
          1152 : Address_next<= 265 ;
          1153 : Address_next<= 132 ;
          1155 : Address_next<= 133 ;
          1156 : Address_next<= 266 ;
          1158 : Address_next<= 267 ;
          1159 : Address_next<= 133 ;
          1160 : Address_next<= 66 ;
          1162 : Address_next<= 67 ;
          1163 : Address_next<= 134 ;
          1164 : Address_next<= 268 ;
          1166 : Address_next<= 269 ;
          1167 : Address_next<= 134 ;
          1169 : Address_next<= 135 ;
          1170 : Address_next<= 270 ;
          1172 : Address_next<= 271 ;
          1173 : Address_next<= 135 ;
          1174 : Address_next<= 67 ;
          1175 : Address_next<= 33 ;
          1176 : Address_next<= 16 ;
          1178 : Address_next<= 17 ;
          1179 : Address_next<= 34 ;
          1180 : Address_next<= 68 ;
          1181 : Address_next<= 136 ;
          1182 : Address_next<= 272 ;
          1184 : Address_next<= 273 ;
          1185 : Address_next<= 136 ;
          1187 : Address_next<= 137 ;
          1188 : Address_next<= 274 ;
          1190 : Address_next<= 275 ;
          1191 : Address_next<= 137 ;
          1192 : Address_next<= 68 ;
          1194 : Address_next<= 69 ;
          1195 : Address_next<= 138 ;
          1196 : Address_next<= 276 ;
          1198 : Address_next<= 277 ;
          1199 : Address_next<= 138 ;
          1201 : Address_next<= 139 ;
          1202 : Address_next<= 278 ;
          1204 : Address_next<= 279 ;
          1205 : Address_next<= 139 ;
          1206 : Address_next<= 69 ;
          1207 : Address_next<= 34 ;
          1209 : Address_next<= 35 ;
          1210 : Address_next<= 70 ;
          1211 : Address_next<= 140 ;
          1212 : Address_next<= 280 ;
          1214 : Address_next<= 281 ;
          1215 : Address_next<= 140 ;
          1217 : Address_next<= 141 ;
          1218 : Address_next<= 282 ;
          1220 : Address_next<= 283 ;
          1221 : Address_next<= 141 ;
          1222 : Address_next<= 70 ;
          1224 : Address_next<= 71 ;
          1225 : Address_next<= 142 ;
          1226 : Address_next<= 284 ;
          1228 : Address_next<= 285 ;
          1229 : Address_next<= 142 ;
          1231 : Address_next<= 143 ;
          1232 : Address_next<= 286 ;
          1234 : Address_next<= 287 ;
          1235 : Address_next<= 143 ;
          1236 : Address_next<= 71 ;
          1237 : Address_next<= 35 ;
          1238 : Address_next<= 17 ;
          1239 : Address_next<= 8 ;
          1242 : Address_next<= 9 ;
          1243 : Address_next<= 18 ;
          1244 : Address_next<= 36 ;
          1245 : Address_next<= 72 ;
          1246 : Address_next<= 144 ;
          1247 : Address_next<= 288 ;
          1249 : Address_next<= 289 ;
          1250 : Address_next<= 144 ;
          1252 : Address_next<= 145 ;
          1253 : Address_next<= 290 ;
          1255 : Address_next<= 291 ;
          1256 : Address_next<= 145 ;
          1257 : Address_next<= 72 ;
          1259 : Address_next<= 73 ;
          1260 : Address_next<= 146 ;
          1261 : Address_next<= 292 ;
          1263 : Address_next<= 293 ;
          1264 : Address_next<= 146 ;
          1266 : Address_next<= 147 ;
          1267 : Address_next<= 294 ;
          1269 : Address_next<= 295 ;
          1270 : Address_next<= 147 ;
          1271 : Address_next<= 73 ;
          1272 : Address_next<= 36 ;
          1274 : Address_next<= 37 ;
          1275 : Address_next<= 74 ;
          1276 : Address_next<= 148 ;
          1277 : Address_next<= 296 ;
          1279 : Address_next<= 297 ;
          1280 : Address_next<= 148 ;
          1282 : Address_next<= 149 ;
          1283 : Address_next<= 298 ;
          1285 : Address_next<= 299 ;
          1286 : Address_next<= 149 ;
          1287 : Address_next<= 74 ;
          1289 : Address_next<= 75 ;
          1290 : Address_next<= 150 ;
          1291 : Address_next<= 300 ;
          1293 : Address_next<= 301 ;
          1294 : Address_next<= 150 ;
          1296 : Address_next<= 151 ;
          1297 : Address_next<= 302 ;
          1299 : Address_next<= 303 ;
          1300 : Address_next<= 151 ;
          1301 : Address_next<= 75 ;
          1302 : Address_next<= 37 ;
          1303 : Address_next<= 18 ;
          1305 : Address_next<= 19 ;
          1306 : Address_next<= 38 ;
          1307 : Address_next<= 76 ;
          1308 : Address_next<= 152 ;
          1309 : Address_next<= 304 ;
          1311 : Address_next<= 305 ;
          1312 : Address_next<= 152 ;
          1314 : Address_next<= 153 ;
          1315 : Address_next<= 306 ;
          1317 : Address_next<= 307 ;
          1318 : Address_next<= 153 ;
          1319 : Address_next<= 76 ;
          1321 : Address_next<= 77 ;
          1322 : Address_next<= 154 ;
          1323 : Address_next<= 308 ;
          1325 : Address_next<= 309 ;
          1326 : Address_next<= 154 ;
          1328 : Address_next<= 155 ;
          1329 : Address_next<= 310 ;
          1331 : Address_next<= 311 ;
          1332 : Address_next<= 155 ;
          1333 : Address_next<= 77 ;
          1334 : Address_next<= 38 ;
          1336 : Address_next<= 39 ;
          1337 : Address_next<= 78 ;
          1338 : Address_next<= 156 ;
          1339 : Address_next<= 312 ;
          1341 : Address_next<= 313 ;
          1342 : Address_next<= 156 ;
          1344 : Address_next<= 157 ;
          1345 : Address_next<= 314 ;
          1347 : Address_next<= 315 ;
          1348 : Address_next<= 157 ;
          1349 : Address_next<= 78 ;
          1351 : Address_next<= 79 ;
          1352 : Address_next<= 158 ;
          1353 : Address_next<= 316 ;
          1355 : Address_next<= 317 ;
          1356 : Address_next<= 158 ;
          1358 : Address_next<= 159 ;
          1359 : Address_next<= 318 ;
          1361 : Address_next<= 319 ;
          1362 : Address_next<= 159 ;
          1363 : Address_next<= 79 ;
          1364 : Address_next<= 39 ;
          1365 : Address_next<= 19 ;
          1366 : Address_next<= 9 ;
          1367 : Address_next<= 4 ;
          1368 : Address_next<= 4 ;
          1373 : Address_next<= 5 ;
          1374 : Address_next<= 5 ;
          1375 : Address_next<= 10 ;
          1376 : Address_next<= 20 ;
          1377 : Address_next<= 40 ;
          1378 : Address_next<= 80 ;
          1379 : Address_next<= 160 ;
          1380 : Address_next<= 320 ;
          1382 : Address_next<= 321 ;
          1383 : Address_next<= 160 ;
          1385 : Address_next<= 161 ;
          1386 : Address_next<= 322 ;
          1388 : Address_next<= 323 ;
          1389 : Address_next<= 161 ;
          1390 : Address_next<= 80 ;
          1392 : Address_next<= 81 ;
          1393 : Address_next<= 162 ;
          1394 : Address_next<= 324 ;
          1396 : Address_next<= 325 ;
          1397 : Address_next<= 162 ;
          1399 : Address_next<= 163 ;
          1400 : Address_next<= 326 ;
          1402 : Address_next<= 327 ;
          1403 : Address_next<= 163 ;
          1404 : Address_next<= 81 ;
          1405 : Address_next<= 40 ;
          1407 : Address_next<= 41 ;
          1408 : Address_next<= 82 ;
          1409 : Address_next<= 164 ;
          1410 : Address_next<= 328 ;
          1412 : Address_next<= 329 ;
          1413 : Address_next<= 164 ;
          1415 : Address_next<= 165 ;
          1416 : Address_next<= 330 ;
          1418 : Address_next<= 331 ;
          1419 : Address_next<= 165 ;
          1420 : Address_next<= 82 ;
          1422 : Address_next<= 83 ;
          1423 : Address_next<= 166 ;
          1424 : Address_next<= 332 ;
          1426 : Address_next<= 333 ;
          1427 : Address_next<= 166 ;
          1429 : Address_next<= 167 ;
          1430 : Address_next<= 334 ;
          1432 : Address_next<= 335 ;
          1433 : Address_next<= 167 ;
          1434 : Address_next<= 83 ;
          1435 : Address_next<= 41 ;
          1436 : Address_next<= 20 ;
          1438 : Address_next<= 21 ;
          1439 : Address_next<= 42 ;
          1440 : Address_next<= 84 ;
          1441 : Address_next<= 168 ;
          1442 : Address_next<= 336 ;
          1444 : Address_next<= 337 ;
          1445 : Address_next<= 168 ;
          1447 : Address_next<= 169 ;
          1448 : Address_next<= 338 ;
          1450 : Address_next<= 339 ;
          1451 : Address_next<= 169 ;
          1452 : Address_next<= 84 ;
          1454 : Address_next<= 85 ;
          1455 : Address_next<= 170 ;
          1456 : Address_next<= 340 ;
          1458 : Address_next<= 341 ;
          1459 : Address_next<= 170 ;
          1461 : Address_next<= 171 ;
          1462 : Address_next<= 342 ;
          1464 : Address_next<= 343 ;
          1465 : Address_next<= 171 ;
          1466 : Address_next<= 85 ;
          1467 : Address_next<= 42 ;
          1469 : Address_next<= 43 ;
          1470 : Address_next<= 86 ;
          1471 : Address_next<= 172 ;
          1472 : Address_next<= 344 ;
          1474 : Address_next<= 345 ;
          1475 : Address_next<= 172 ;
          1477 : Address_next<= 173 ;
          1478 : Address_next<= 346 ;
          1480 : Address_next<= 347 ;
          1481 : Address_next<= 173 ;
          1482 : Address_next<= 86 ;
          1484 : Address_next<= 87 ;
          1485 : Address_next<= 174 ;
          1486 : Address_next<= 348 ;
          1488 : Address_next<= 349 ;
          1489 : Address_next<= 174 ;
          1491 : Address_next<= 175 ;
          1492 : Address_next<= 350 ;
          1494 : Address_next<= 351 ;
          1495 : Address_next<= 175 ;
          1496 : Address_next<= 87 ;
          1497 : Address_next<= 43 ;
          1498 : Address_next<= 21 ;
          1499 : Address_next<= 10 ;
          1502 : Address_next<= 11 ;
          1503 : Address_next<= 22 ;
          1504 : Address_next<= 44 ;
          1505 : Address_next<= 88 ;
          1506 : Address_next<= 176 ;
          1507 : Address_next<= 352 ;
          1509 : Address_next<= 353 ;
          1510 : Address_next<= 176 ;
          1512 : Address_next<= 177 ;
          1513 : Address_next<= 354 ;
          1515 : Address_next<= 355 ;
          1516 : Address_next<= 177 ;
          1517 : Address_next<= 88 ;
          1519 : Address_next<= 89 ;
          1520 : Address_next<= 178 ;
          1521 : Address_next<= 356 ;
          1523 : Address_next<= 357 ;
          1524 : Address_next<= 178 ;
          1526 : Address_next<= 179 ;
          1527 : Address_next<= 358 ;
          1529 : Address_next<= 359 ;
          1530 : Address_next<= 179 ;
          1531 : Address_next<= 89 ;
          1532 : Address_next<= 44 ;
          1534 : Address_next<= 45 ;
          1535 : Address_next<= 90 ;
          1536 : Address_next<= 180 ;
          1537 : Address_next<= 360 ;
          1539 : Address_next<= 361 ;
          1540 : Address_next<= 180 ;
          1542 : Address_next<= 181 ;
          1543 : Address_next<= 362 ;
          1545 : Address_next<= 363 ;
          1546 : Address_next<= 181 ;
          1547 : Address_next<= 90 ;
          1549 : Address_next<= 91 ;
          1550 : Address_next<= 182 ;
          1551 : Address_next<= 364 ;
          1553 : Address_next<= 365 ;
          1554 : Address_next<= 182 ;
          1556 : Address_next<= 183 ;
          1557 : Address_next<= 366 ;
          1559 : Address_next<= 367 ;
          1560 : Address_next<= 183 ;
          1561 : Address_next<= 91 ;
          1562 : Address_next<= 45 ;
          1563 : Address_next<= 22 ;
          1565 : Address_next<= 23 ;
          1566 : Address_next<= 46 ;
          1567 : Address_next<= 92 ;
          1568 : Address_next<= 184 ;
          1569 : Address_next<= 368 ;
          1571 : Address_next<= 369 ;
          1572 : Address_next<= 184 ;
          1574 : Address_next<= 185 ;
          1575 : Address_next<= 370 ;
          1577 : Address_next<= 371 ;
          1578 : Address_next<= 185 ;
          1579 : Address_next<= 92 ;
          1581 : Address_next<= 93 ;
          1582 : Address_next<= 186 ;
          1583 : Address_next<= 372 ;
          1585 : Address_next<= 373 ;
          1586 : Address_next<= 186 ;
          1588 : Address_next<= 187 ;
          1589 : Address_next<= 374 ;
          1591 : Address_next<= 375 ;
          1592 : Address_next<= 187 ;
          1593 : Address_next<= 93 ;
          1594 : Address_next<= 46 ;
          1596 : Address_next<= 47 ;
          1597 : Address_next<= 94 ;
          1598 : Address_next<= 188 ;
          1599 : Address_next<= 376 ;
          1601 : Address_next<= 377 ;
          1602 : Address_next<= 188 ;
          1604 : Address_next<= 189 ;
          1605 : Address_next<= 378 ;
          1607 : Address_next<= 379 ;
          1608 : Address_next<= 189 ;
          1609 : Address_next<= 94 ;
          1611 : Address_next<= 95 ;
          1612 : Address_next<= 190 ;
          1613 : Address_next<= 380 ;
          1615 : Address_next<= 381 ;
          1616 : Address_next<= 190 ;
          1618 : Address_next<= 191 ;
          1619 : Address_next<= 382 ;
          1621 : Address_next<= 383 ;
          1622 : Address_next<= 191 ;
          1623 : Address_next<= 95 ;
          1624 : Address_next<= 47 ;
          1625 : Address_next<= 23 ;
          1626 : Address_next<= 11 ;
          1627 : Address_next<= 5 ;
          1628 : Address_next<= 5 ;
          1629 : Address_next<= 2 ;
          1630 : Address_next<= 2 ;
          1631 : Address_next<= 2 ;
          1632 : Address_next<= 2 ;
          1641 : Address_next<= 3 ;
          1642 : Address_next<= 3 ;
          1643 : Address_next<= 3 ;
          1644 : Address_next<= 3 ;
          1645 : Address_next<= 6 ;
          1646 : Address_next<= 6 ;
          1647 : Address_next<= 12 ;
          1648 : Address_next<= 24 ;
          1649 : Address_next<= 48 ;
          1650 : Address_next<= 96 ;
          1651 : Address_next<= 192 ;
          1652 : Address_next<= 384 ;
          1654 : Address_next<= 385 ;
          1655 : Address_next<= 192 ;
          1657 : Address_next<= 193 ;
          1658 : Address_next<= 386 ;
          1660 : Address_next<= 387 ;
          1661 : Address_next<= 193 ;
          1662 : Address_next<= 96 ;
          1664 : Address_next<= 97 ;
          1665 : Address_next<= 194 ;
          1666 : Address_next<= 388 ;
          1668 : Address_next<= 389 ;
          1669 : Address_next<= 194 ;
          1671 : Address_next<= 195 ;
          1672 : Address_next<= 390 ;
          1674 : Address_next<= 391 ;
          1675 : Address_next<= 195 ;
          1676 : Address_next<= 97 ;
          1677 : Address_next<= 48 ;
          1679 : Address_next<= 49 ;
          1680 : Address_next<= 98 ;
          1681 : Address_next<= 196 ;
          1682 : Address_next<= 392 ;
          1684 : Address_next<= 393 ;
          1685 : Address_next<= 196 ;
          1687 : Address_next<= 197 ;
          1688 : Address_next<= 394 ;
          1690 : Address_next<= 395 ;
          1691 : Address_next<= 197 ;
          1692 : Address_next<= 98 ;
          1694 : Address_next<= 99 ;
          1695 : Address_next<= 198 ;
          1696 : Address_next<= 396 ;
          1698 : Address_next<= 397 ;
          1699 : Address_next<= 198 ;
          1701 : Address_next<= 199 ;
          1702 : Address_next<= 398 ;
          1704 : Address_next<= 399 ;
          1705 : Address_next<= 199 ;
          1706 : Address_next<= 99 ;
          1707 : Address_next<= 49 ;
          1708 : Address_next<= 24 ;
          1710 : Address_next<= 25 ;
          1711 : Address_next<= 50 ;
          1712 : Address_next<= 100 ;
          1713 : Address_next<= 200 ;
          1714 : Address_next<= 400 ;
          1716 : Address_next<= 401 ;
          1717 : Address_next<= 200 ;
          1719 : Address_next<= 201 ;
          1720 : Address_next<= 402 ;
          1722 : Address_next<= 403 ;
          1723 : Address_next<= 201 ;
          1724 : Address_next<= 100 ;
          1726 : Address_next<= 101 ;
          1727 : Address_next<= 202 ;
          1728 : Address_next<= 404 ;
          1730 : Address_next<= 405 ;
          1731 : Address_next<= 202 ;
          1733 : Address_next<= 203 ;
          1734 : Address_next<= 406 ;
          1736 : Address_next<= 407 ;
          1737 : Address_next<= 203 ;
          1738 : Address_next<= 101 ;
          1739 : Address_next<= 50 ;
          1741 : Address_next<= 51 ;
          1742 : Address_next<= 102 ;
          1743 : Address_next<= 204 ;
          1744 : Address_next<= 408 ;
          1746 : Address_next<= 409 ;
          1747 : Address_next<= 204 ;
          1749 : Address_next<= 205 ;
          1750 : Address_next<= 410 ;
          1752 : Address_next<= 411 ;
          1753 : Address_next<= 205 ;
          1754 : Address_next<= 102 ;
          1756 : Address_next<= 103 ;
          1757 : Address_next<= 206 ;
          1758 : Address_next<= 412 ;
          1760 : Address_next<= 413 ;
          1761 : Address_next<= 206 ;
          1763 : Address_next<= 207 ;
          1764 : Address_next<= 414 ;
          1766 : Address_next<= 415 ;
          1767 : Address_next<= 207 ;
          1768 : Address_next<= 103 ;
          1769 : Address_next<= 51 ;
          1770 : Address_next<= 25 ;
          1771 : Address_next<= 12 ;
          1774 : Address_next<= 13 ;
          1775 : Address_next<= 26 ;
          1776 : Address_next<= 52 ;
          1777 : Address_next<= 104 ;
          1778 : Address_next<= 208 ;
          1779 : Address_next<= 416 ;
          1781 : Address_next<= 417 ;
          1782 : Address_next<= 208 ;
          1784 : Address_next<= 209 ;
          1785 : Address_next<= 418 ;
          1787 : Address_next<= 419 ;
          1788 : Address_next<= 209 ;
          1789 : Address_next<= 104 ;
          1791 : Address_next<= 105 ;
          1792 : Address_next<= 210 ;
          1793 : Address_next<= 420 ;
          1795 : Address_next<= 421 ;
          1796 : Address_next<= 210 ;
          1798 : Address_next<= 211 ;
          1799 : Address_next<= 422 ;
          1801 : Address_next<= 423 ;
          1802 : Address_next<= 211 ;
          1803 : Address_next<= 105 ;
          1804 : Address_next<= 52 ;
          1806 : Address_next<= 53 ;
          1807 : Address_next<= 106 ;
          1808 : Address_next<= 212 ;
          1809 : Address_next<= 424 ;
          1811 : Address_next<= 425 ;
          1812 : Address_next<= 212 ;
          1814 : Address_next<= 213 ;
          1815 : Address_next<= 426 ;
          1817 : Address_next<= 427 ;
          1818 : Address_next<= 213 ;
          1819 : Address_next<= 106 ;
          1821 : Address_next<= 107 ;
          1822 : Address_next<= 214 ;
          1823 : Address_next<= 428 ;
          1825 : Address_next<= 429 ;
          1826 : Address_next<= 214 ;
          1828 : Address_next<= 215 ;
          1829 : Address_next<= 430 ;
          1831 : Address_next<= 431 ;
          1832 : Address_next<= 215 ;
          1833 : Address_next<= 107 ;
          1834 : Address_next<= 53 ;
          1835 : Address_next<= 26 ;
          1837 : Address_next<= 27 ;
          1838 : Address_next<= 54 ;
          1839 : Address_next<= 108 ;
          1840 : Address_next<= 216 ;
          1841 : Address_next<= 432 ;
          1843 : Address_next<= 433 ;
          1844 : Address_next<= 216 ;
          1846 : Address_next<= 217 ;
          1847 : Address_next<= 434 ;
          1849 : Address_next<= 435 ;
          1850 : Address_next<= 217 ;
          1851 : Address_next<= 108 ;
          1853 : Address_next<= 109 ;
          1854 : Address_next<= 218 ;
          1855 : Address_next<= 436 ;
          1857 : Address_next<= 437 ;
          1858 : Address_next<= 218 ;
          1860 : Address_next<= 219 ;
          1861 : Address_next<= 438 ;
          1863 : Address_next<= 439 ;
          1864 : Address_next<= 219 ;
          1865 : Address_next<= 109 ;
          1866 : Address_next<= 54 ;
          1868 : Address_next<= 55 ;
          1869 : Address_next<= 110 ;
          1870 : Address_next<= 220 ;
          1871 : Address_next<= 440 ;
          1873 : Address_next<= 441 ;
          1874 : Address_next<= 220 ;
          1876 : Address_next<= 221 ;
          1877 : Address_next<= 442 ;
          1879 : Address_next<= 443 ;
          1880 : Address_next<= 221 ;
          1881 : Address_next<= 110 ;
          1883 : Address_next<= 111 ;
          1884 : Address_next<= 222 ;
          1885 : Address_next<= 444 ;
          1887 : Address_next<= 445 ;
          1888 : Address_next<= 222 ;
          1890 : Address_next<= 223 ;
          1891 : Address_next<= 446 ;
          1893 : Address_next<= 447 ;
          1894 : Address_next<= 223 ;
          1895 : Address_next<= 111 ;
          1896 : Address_next<= 55 ;
          1897 : Address_next<= 27 ;
          1898 : Address_next<= 13 ;
          1899 : Address_next<= 6 ;
          1900 : Address_next<= 6 ;
          1905 : Address_next<= 7 ;
          1906 : Address_next<= 7 ;
          1907 : Address_next<= 14 ;
          1908 : Address_next<= 28 ;
          1909 : Address_next<= 56 ;
          1910 : Address_next<= 112 ;
          1911 : Address_next<= 224 ;
          1912 : Address_next<= 448 ;
          1914 : Address_next<= 449 ;
          1915 : Address_next<= 224 ;
          1917 : Address_next<= 225 ;
          1918 : Address_next<= 450 ;
          1920 : Address_next<= 451 ;
          1921 : Address_next<= 225 ;
          1922 : Address_next<= 112 ;
          1924 : Address_next<= 113 ;
          1925 : Address_next<= 226 ;
          1926 : Address_next<= 452 ;
          1928 : Address_next<= 453 ;
          1929 : Address_next<= 226 ;
          1931 : Address_next<= 227 ;
          1932 : Address_next<= 454 ;
          1934 : Address_next<= 455 ;
          1935 : Address_next<= 227 ;
          1936 : Address_next<= 113 ;
          1937 : Address_next<= 56 ;
          1939 : Address_next<= 57 ;
          1940 : Address_next<= 114 ;
          1941 : Address_next<= 228 ;
          1942 : Address_next<= 456 ;
          1944 : Address_next<= 457 ;
          1945 : Address_next<= 228 ;
          1947 : Address_next<= 229 ;
          1948 : Address_next<= 458 ;
          1950 : Address_next<= 459 ;
          1951 : Address_next<= 229 ;
          1952 : Address_next<= 114 ;
          1954 : Address_next<= 115 ;
          1955 : Address_next<= 230 ;
          1956 : Address_next<= 460 ;
          1958 : Address_next<= 461 ;
          1959 : Address_next<= 230 ;
          1961 : Address_next<= 231 ;
          1962 : Address_next<= 462 ;
          1964 : Address_next<= 463 ;
          1965 : Address_next<= 231 ;
          1966 : Address_next<= 115 ;
          1967 : Address_next<= 57 ;
          1968 : Address_next<= 28 ;
          1970 : Address_next<= 29 ;
          1971 : Address_next<= 58 ;
          1972 : Address_next<= 116 ;
          1973 : Address_next<= 232 ;
          1974 : Address_next<= 464 ;
          1976 : Address_next<= 465 ;
          1977 : Address_next<= 232 ;
          1979 : Address_next<= 233 ;
          1980 : Address_next<= 466 ;
          1982 : Address_next<= 467 ;
          1983 : Address_next<= 233 ;
          1984 : Address_next<= 116 ;
          1986 : Address_next<= 117 ;
          1987 : Address_next<= 234 ;
          1988 : Address_next<= 468 ;
          1990 : Address_next<= 469 ;
          1991 : Address_next<= 234 ;
          1993 : Address_next<= 235 ;
          1994 : Address_next<= 470 ;
          1996 : Address_next<= 471 ;
          1997 : Address_next<= 235 ;
          1998 : Address_next<= 117 ;
          1999 : Address_next<= 58 ;
          2001 : Address_next<= 59 ;
          2002 : Address_next<= 118 ;
          2003 : Address_next<= 236 ;
          2004 : Address_next<= 472 ;
          2006 : Address_next<= 473 ;
          2007 : Address_next<= 236 ;
          2009 : Address_next<= 237 ;
          2010 : Address_next<= 474 ;
          2012 : Address_next<= 475 ;
          2013 : Address_next<= 237 ;
          2014 : Address_next<= 118 ;
          2016 : Address_next<= 119 ;
          2017 : Address_next<= 238 ;
          2018 : Address_next<= 476 ;
          2020 : Address_next<= 477 ;
          2021 : Address_next<= 238 ;
          2023 : Address_next<= 239 ;
          2024 : Address_next<= 478 ;
          2026 : Address_next<= 479 ;
          2027 : Address_next<= 239 ;
          2028 : Address_next<= 119 ;
          2029 : Address_next<= 59 ;
          2030 : Address_next<= 29 ;
          2031 : Address_next<= 14 ;
          2034 : Address_next<= 15 ;
          2035 : Address_next<= 30 ;
          2036 : Address_next<= 60 ;
          2037 : Address_next<= 120 ;
          2038 : Address_next<= 240 ;
          2039 : Address_next<= 480 ;
          2041 : Address_next<= 481 ;
          2042 : Address_next<= 240 ;
          2044 : Address_next<= 241 ;
          2045 : Address_next<= 482 ;
          2047 : Address_next<= 483 ;
          2048 : Address_next<= 241 ;
          2049 : Address_next<= 120 ;
          2051 : Address_next<= 121 ;
          2052 : Address_next<= 242 ;
          2053 : Address_next<= 484 ;
          2055 : Address_next<= 485 ;
          2056 : Address_next<= 242 ;
          2058 : Address_next<= 243 ;
          2059 : Address_next<= 486 ;
          2061 : Address_next<= 487 ;
          2062 : Address_next<= 243 ;
          2063 : Address_next<= 121 ;
          2064 : Address_next<= 60 ;
          2066 : Address_next<= 61 ;
          2067 : Address_next<= 122 ;
          2068 : Address_next<= 244 ;
          2069 : Address_next<= 488 ;
          2071 : Address_next<= 489 ;
          2072 : Address_next<= 244 ;
          2074 : Address_next<= 245 ;
          2075 : Address_next<= 490 ;
          2077 : Address_next<= 491 ;
          2078 : Address_next<= 245 ;
          2079 : Address_next<= 122 ;
          2081 : Address_next<= 123 ;
          2082 : Address_next<= 246 ;
          2083 : Address_next<= 492 ;
          2085 : Address_next<= 493 ;
          2086 : Address_next<= 246 ;
          2088 : Address_next<= 247 ;
          2089 : Address_next<= 494 ;
          2091 : Address_next<= 495 ;
          2092 : Address_next<= 247 ;
          2093 : Address_next<= 123 ;
          2094 : Address_next<= 61 ;
          2095 : Address_next<= 30 ;
          2097 : Address_next<= 31 ;
          2098 : Address_next<= 62 ;
          2099 : Address_next<= 124 ;
          2100 : Address_next<= 248 ;
          2101 : Address_next<= 496 ;
          2103 : Address_next<= 497 ;
          2104 : Address_next<= 248 ;
          2106 : Address_next<= 249 ;
          2107 : Address_next<= 498 ;
          2109 : Address_next<= 499 ;
          2110 : Address_next<= 249 ;
          2111 : Address_next<= 124 ;
          2113 : Address_next<= 125 ;
          2114 : Address_next<= 250 ;
          2115 : Address_next<= 500 ;
          2117 : Address_next<= 501 ;
          2118 : Address_next<= 250 ;
          2120 : Address_next<= 251 ;
          2121 : Address_next<= 502 ;
          2123 : Address_next<= 503 ;
          2124 : Address_next<= 251 ;
          2125 : Address_next<= 125 ;
          2126 : Address_next<= 62 ;
          2128 : Address_next<= 63 ;
          2129 : Address_next<= 126 ;
          2130 : Address_next<= 252 ;
          2131 : Address_next<= 504 ;
          2133 : Address_next<= 505 ;
          2134 : Address_next<= 252 ;
          2136 : Address_next<= 253 ;
          2137 : Address_next<= 506 ;
          2139 : Address_next<= 507 ;
          2140 : Address_next<= 253 ;
          2141 : Address_next<= 126 ;
          2143 : Address_next<= 127 ;
          2144 : Address_next<= 254 ;
          2145 : Address_next<= 508 ;
          2147 : Address_next<= 509 ;
          2148 : Address_next<= 254 ;
          2150 : Address_next<= 255 ;
          2151 : Address_next<= 510 ;
          2153 : Address_next<= 511 ;
          2154 : Address_next<= 255 ;
          2155 : Address_next<= 127 ;
          2156 : Address_next<= 63 ;
          2157 : Address_next<= 31 ;
          2158 : Address_next<= 15 ;
          2159 : Address_next<= 7 ;
          2160 : Address_next<= 7 ;
          2161 : Address_next<= 3 ;
          2162 : Address_next<= 3 ;
          2163 : Address_next<= 3 ;
          2164 : Address_next<= 3 ;
          2165 : Address_next<= 1 ;
          2166 : Address_next<= 1 ;
          2167 : Address_next<= 1 ;
          2168 : Address_next<= 1 ;
          2169 : Address_next<= 1 ;
          2170 : Address_next<= 1 ;
          2171 : Address_next<= 1 ;
          2172 : Address_next<= 1 ;
       endcase









      end
      else begin
           L_Nv_next                     <=1024;
           L_opcode_next <= TYPE1;
           L_part_count_next <= 0;
           Address_next <= 0;
      end
end
end
endmodule


