module frozen_rom 
(input [12:0] in_bit_index, input en, output frozen1,output frozen2, input clk);
wire [12:0] in_bit_index2;
 assign in_bit_index2 = in_bit_index + 1 ;
reg out, out2;
 assign frozen1 = out;
 assign frozen2 = out2;
always @(posedge clk) begin
if (en) begin
case(in_bit_index)
  0 :out<= 0 ;
  1 :out<= 0 ;
  2 :out<= 0 ;
  3 :out<= 0 ;
  4 :out<= 0 ;
  5 :out<= 0 ;
  6 :out<= 0 ;
  7 :out<= 0 ;
  8 :out<= 0 ;
  9 :out<= 0 ;
  10 :out<= 0 ;
  11 :out<= 0 ;
  12 :out<= 0 ;
  13 :out<= 0 ;
  14 :out<= 0 ;
  15 :out<= 0 ;
  16 :out<= 0 ;
  17 :out<= 0 ;
  18 :out<= 0 ;
  19 :out<= 0 ;
  20 :out<= 0 ;
  21 :out<= 0 ;
  22 :out<= 0 ;
  23 :out<= 0 ;
  24 :out<= 0 ;
  25 :out<= 0 ;
  26 :out<= 0 ;
  27 :out<= 0 ;
  28 :out<= 0 ;
  29 :out<= 0 ;
  30 :out<= 0 ;
  31 :out<= 0 ;
  32 :out<= 0 ;
  33 :out<= 0 ;
  34 :out<= 0 ;
  35 :out<= 0 ;
  36 :out<= 0 ;
  37 :out<= 0 ;
  38 :out<= 0 ;
  39 :out<= 0 ;
  40 :out<= 0 ;
  41 :out<= 0 ;
  42 :out<= 0 ;
  43 :out<= 0 ;
  44 :out<= 0 ;
  45 :out<= 0 ;
  46 :out<= 0 ;
  47 :out<= 0 ;
  48 :out<= 0 ;
  49 :out<= 0 ;
  50 :out<= 0 ;
  51 :out<= 0 ;
  52 :out<= 0 ;
  53 :out<= 0 ;
  54 :out<= 0 ;
  55 :out<= 0 ;
  56 :out<= 0 ;
  57 :out<= 0 ;
  58 :out<= 0 ;
  59 :out<= 0 ;
  60 :out<= 0 ;
  61 :out<= 0 ;
  62 :out<= 0 ;
  63 :out<= 0 ;
  64 :out<= 0 ;
  65 :out<= 0 ;
  66 :out<= 0 ;
  67 :out<= 0 ;
  68 :out<= 0 ;
  69 :out<= 0 ;
  70 :out<= 0 ;
  71 :out<= 0 ;
  72 :out<= 0 ;
  73 :out<= 0 ;
  74 :out<= 0 ;
  75 :out<= 0 ;
  76 :out<= 0 ;
  77 :out<= 0 ;
  78 :out<= 0 ;
  79 :out<= 0 ;
  80 :out<= 0 ;
  81 :out<= 0 ;
  82 :out<= 0 ;
  83 :out<= 0 ;
  84 :out<= 0 ;
  85 :out<= 0 ;
  86 :out<= 0 ;
  87 :out<= 0 ;
  88 :out<= 0 ;
  89 :out<= 0 ;
  90 :out<= 0 ;
  91 :out<= 0 ;
  92 :out<= 0 ;
  93 :out<= 0 ;
  94 :out<= 0 ;
  95 :out<= 0 ;
  96 :out<= 0 ;
  97 :out<= 0 ;
  98 :out<= 0 ;
  99 :out<= 0 ;
  100 :out<= 0 ;
  101 :out<= 0 ;
  102 :out<= 0 ;
  103 :out<= 0 ;
  104 :out<= 0 ;
  105 :out<= 0 ;
  106 :out<= 0 ;
  107 :out<= 0 ;
  108 :out<= 0 ;
  109 :out<= 0 ;
  110 :out<= 0 ;
  111 :out<= 0 ;
  112 :out<= 0 ;
  113 :out<= 0 ;
  114 :out<= 0 ;
  115 :out<= 0 ;
  116 :out<= 0 ;
  117 :out<= 0 ;
  118 :out<= 0 ;
  119 :out<= 0 ;
  120 :out<= 0 ;
  121 :out<= 0 ;
  122 :out<= 0 ;
  123 :out<= 0 ;
  124 :out<= 0 ;
  125 :out<= 0 ;
  126 :out<= 0 ;
  127 :out<= 0 ;
  128 :out<= 0 ;
  129 :out<= 0 ;
  130 :out<= 0 ;
  131 :out<= 0 ;
  132 :out<= 0 ;
  133 :out<= 0 ;
  134 :out<= 0 ;
  135 :out<= 0 ;
  136 :out<= 0 ;
  137 :out<= 0 ;
  138 :out<= 0 ;
  139 :out<= 0 ;
  140 :out<= 0 ;
  141 :out<= 0 ;
  142 :out<= 0 ;
  143 :out<= 0 ;
  144 :out<= 0 ;
  145 :out<= 0 ;
  146 :out<= 0 ;
  147 :out<= 0 ;
  148 :out<= 0 ;
  149 :out<= 0 ;
  150 :out<= 0 ;
  151 :out<= 0 ;
  152 :out<= 0 ;
  153 :out<= 0 ;
  154 :out<= 0 ;
  155 :out<= 0 ;
  156 :out<= 0 ;
  157 :out<= 0 ;
  158 :out<= 0 ;
  159 :out<= 0 ;
  160 :out<= 0 ;
  161 :out<= 0 ;
  162 :out<= 0 ;
  163 :out<= 0 ;
  164 :out<= 0 ;
  165 :out<= 0 ;
  166 :out<= 0 ;
  167 :out<= 0 ;
  168 :out<= 0 ;
  169 :out<= 0 ;
  170 :out<= 0 ;
  171 :out<= 0 ;
  172 :out<= 0 ;
  173 :out<= 0 ;
  174 :out<= 0 ;
  175 :out<= 0 ;
  176 :out<= 0 ;
  177 :out<= 0 ;
  178 :out<= 0 ;
  179 :out<= 0 ;
  180 :out<= 0 ;
  181 :out<= 0 ;
  182 :out<= 0 ;
  183 :out<= 0 ;
  184 :out<= 0 ;
  185 :out<= 0 ;
  186 :out<= 0 ;
  187 :out<= 0 ;
  188 :out<= 0 ;
  189 :out<= 0 ;
  190 :out<= 0 ;
  191 :out<= 1 ;
  192 :out<= 0 ;
  193 :out<= 0 ;
  194 :out<= 0 ;
  195 :out<= 0 ;
  196 :out<= 0 ;
  197 :out<= 0 ;
  198 :out<= 0 ;
  199 :out<= 0 ;
  200 :out<= 0 ;
  201 :out<= 0 ;
  202 :out<= 0 ;
  203 :out<= 0 ;
  204 :out<= 0 ;
  205 :out<= 0 ;
  206 :out<= 0 ;
  207 :out<= 0 ;
  208 :out<= 0 ;
  209 :out<= 0 ;
  210 :out<= 0 ;
  211 :out<= 0 ;
  212 :out<= 0 ;
  213 :out<= 0 ;
  214 :out<= 0 ;
  215 :out<= 0 ;
  216 :out<= 0 ;
  217 :out<= 0 ;
  218 :out<= 0 ;
  219 :out<= 0 ;
  220 :out<= 0 ;
  221 :out<= 0 ;
  222 :out<= 0 ;
  223 :out<= 1 ;
  224 :out<= 0 ;
  225 :out<= 0 ;
  226 :out<= 0 ;
  227 :out<= 0 ;
  228 :out<= 0 ;
  229 :out<= 0 ;
  230 :out<= 0 ;
  231 :out<= 0 ;
  232 :out<= 0 ;
  233 :out<= 0 ;
  234 :out<= 0 ;
  235 :out<= 1 ;
  236 :out<= 0 ;
  237 :out<= 1 ;
  238 :out<= 1 ;
  239 :out<= 1 ;
  240 :out<= 0 ;
  241 :out<= 0 ;
  242 :out<= 0 ;
  243 :out<= 1 ;
  244 :out<= 0 ;
  245 :out<= 1 ;
  246 :out<= 1 ;
  247 :out<= 1 ;
  248 :out<= 0 ;
  249 :out<= 1 ;
  250 :out<= 1 ;
  251 :out<= 1 ;
  252 :out<= 1 ;
  253 :out<= 1 ;
  254 :out<= 1 ;
  255 :out<= 1 ;
  256 :out<= 0 ;
  257 :out<= 0 ;
  258 :out<= 0 ;
  259 :out<= 0 ;
  260 :out<= 0 ;
  261 :out<= 0 ;
  262 :out<= 0 ;
  263 :out<= 0 ;
  264 :out<= 0 ;
  265 :out<= 0 ;
  266 :out<= 0 ;
  267 :out<= 0 ;
  268 :out<= 0 ;
  269 :out<= 0 ;
  270 :out<= 0 ;
  271 :out<= 0 ;
  272 :out<= 0 ;
  273 :out<= 0 ;
  274 :out<= 0 ;
  275 :out<= 0 ;
  276 :out<= 0 ;
  277 :out<= 0 ;
  278 :out<= 0 ;
  279 :out<= 0 ;
  280 :out<= 0 ;
  281 :out<= 0 ;
  282 :out<= 0 ;
  283 :out<= 0 ;
  284 :out<= 0 ;
  285 :out<= 0 ;
  286 :out<= 0 ;
  287 :out<= 0 ;
  288 :out<= 0 ;
  289 :out<= 0 ;
  290 :out<= 0 ;
  291 :out<= 0 ;
  292 :out<= 0 ;
  293 :out<= 0 ;
  294 :out<= 0 ;
  295 :out<= 0 ;
  296 :out<= 0 ;
  297 :out<= 0 ;
  298 :out<= 0 ;
  299 :out<= 0 ;
  300 :out<= 0 ;
  301 :out<= 0 ;
  302 :out<= 0 ;
  303 :out<= 0 ;
  304 :out<= 0 ;
  305 :out<= 0 ;
  306 :out<= 0 ;
  307 :out<= 0 ;
  308 :out<= 0 ;
  309 :out<= 0 ;
  310 :out<= 0 ;
  311 :out<= 0 ;
  312 :out<= 0 ;
  313 :out<= 0 ;
  314 :out<= 0 ;
  315 :out<= 1 ;
  316 :out<= 0 ;
  317 :out<= 1 ;
  318 :out<= 1 ;
  319 :out<= 1 ;
  320 :out<= 0 ;
  321 :out<= 0 ;
  322 :out<= 0 ;
  323 :out<= 0 ;
  324 :out<= 0 ;
  325 :out<= 0 ;
  326 :out<= 0 ;
  327 :out<= 0 ;
  328 :out<= 0 ;
  329 :out<= 0 ;
  330 :out<= 0 ;
  331 :out<= 0 ;
  332 :out<= 0 ;
  333 :out<= 0 ;
  334 :out<= 0 ;
  335 :out<= 0 ;
  336 :out<= 0 ;
  337 :out<= 0 ;
  338 :out<= 0 ;
  339 :out<= 0 ;
  340 :out<= 0 ;
  341 :out<= 0 ;
  342 :out<= 0 ;
  343 :out<= 1 ;
  344 :out<= 0 ;
  345 :out<= 0 ;
  346 :out<= 0 ;
  347 :out<= 1 ;
  348 :out<= 0 ;
  349 :out<= 1 ;
  350 :out<= 1 ;
  351 :out<= 1 ;
  352 :out<= 0 ;
  353 :out<= 0 ;
  354 :out<= 0 ;
  355 :out<= 0 ;
  356 :out<= 0 ;
  357 :out<= 0 ;
  358 :out<= 0 ;
  359 :out<= 1 ;
  360 :out<= 0 ;
  361 :out<= 0 ;
  362 :out<= 0 ;
  363 :out<= 1 ;
  364 :out<= 0 ;
  365 :out<= 1 ;
  366 :out<= 1 ;
  367 :out<= 1 ;
  368 :out<= 0 ;
  369 :out<= 0 ;
  370 :out<= 1 ;
  371 :out<= 1 ;
  372 :out<= 1 ;
  373 :out<= 1 ;
  374 :out<= 1 ;
  375 :out<= 1 ;
  376 :out<= 1 ;
  377 :out<= 1 ;
  378 :out<= 1 ;
  379 :out<= 1 ;
  380 :out<= 1 ;
  381 :out<= 1 ;
  382 :out<= 1 ;
  383 :out<= 1 ;
  384 :out<= 0 ;
  385 :out<= 0 ;
  386 :out<= 0 ;
  387 :out<= 0 ;
  388 :out<= 0 ;
  389 :out<= 0 ;
  390 :out<= 0 ;
  391 :out<= 0 ;
  392 :out<= 0 ;
  393 :out<= 0 ;
  394 :out<= 0 ;
  395 :out<= 0 ;
  396 :out<= 0 ;
  397 :out<= 0 ;
  398 :out<= 0 ;
  399 :out<= 1 ;
  400 :out<= 0 ;
  401 :out<= 0 ;
  402 :out<= 0 ;
  403 :out<= 0 ;
  404 :out<= 0 ;
  405 :out<= 0 ;
  406 :out<= 0 ;
  407 :out<= 1 ;
  408 :out<= 0 ;
  409 :out<= 0 ;
  410 :out<= 1 ;
  411 :out<= 1 ;
  412 :out<= 1 ;
  413 :out<= 1 ;
  414 :out<= 1 ;
  415 :out<= 1 ;
  416 :out<= 0 ;
  417 :out<= 0 ;
  418 :out<= 0 ;
  419 :out<= 0 ;
  420 :out<= 0 ;
  421 :out<= 1 ;
  422 :out<= 1 ;
  423 :out<= 1 ;
  424 :out<= 0 ;
  425 :out<= 1 ;
  426 :out<= 1 ;
  427 :out<= 1 ;
  428 :out<= 1 ;
  429 :out<= 1 ;
  430 :out<= 1 ;
  431 :out<= 1 ;
  432 :out<= 0 ;
  433 :out<= 1 ;
  434 :out<= 1 ;
  435 :out<= 1 ;
  436 :out<= 1 ;
  437 :out<= 1 ;
  438 :out<= 1 ;
  439 :out<= 1 ;
  440 :out<= 1 ;
  441 :out<= 1 ;
  442 :out<= 1 ;
  443 :out<= 1 ;
  444 :out<= 1 ;
  445 :out<= 1 ;
  446 :out<= 1 ;
  447 :out<= 1 ;
  448 :out<= 0 ;
  449 :out<= 0 ;
  450 :out<= 0 ;
  451 :out<= 1 ;
  452 :out<= 0 ;
  453 :out<= 1 ;
  454 :out<= 1 ;
  455 :out<= 1 ;
  456 :out<= 0 ;
  457 :out<= 1 ;
  458 :out<= 1 ;
  459 :out<= 1 ;
  460 :out<= 1 ;
  461 :out<= 1 ;
  462 :out<= 1 ;
  463 :out<= 1 ;
  464 :out<= 0 ;
  465 :out<= 1 ;
  466 :out<= 1 ;
  467 :out<= 1 ;
  468 :out<= 1 ;
  469 :out<= 1 ;
  470 :out<= 1 ;
  471 :out<= 1 ;
  472 :out<= 1 ;
  473 :out<= 1 ;
  474 :out<= 1 ;
  475 :out<= 1 ;
  476 :out<= 1 ;
  477 :out<= 1 ;
  478 :out<= 1 ;
  479 :out<= 1 ;
  480 :out<= 0 ;
  481 :out<= 1 ;
  482 :out<= 1 ;
  483 :out<= 1 ;
  484 :out<= 1 ;
  485 :out<= 1 ;
  486 :out<= 1 ;
  487 :out<= 1 ;
  488 :out<= 1 ;
  489 :out<= 1 ;
  490 :out<= 1 ;
  491 :out<= 1 ;
  492 :out<= 1 ;
  493 :out<= 1 ;
  494 :out<= 1 ;
  495 :out<= 1 ;
  496 :out<= 1 ;
  497 :out<= 1 ;
  498 :out<= 1 ;
  499 :out<= 1 ;
  500 :out<= 1 ;
  501 :out<= 1 ;
  502 :out<= 1 ;
  503 :out<= 1 ;
  504 :out<= 1 ;
  505 :out<= 1 ;
  506 :out<= 1 ;
  507 :out<= 1 ;
  508 :out<= 1 ;
  509 :out<= 1 ;
  510 :out<= 1 ;
  511 :out<= 1 ;
  512 :out<= 0 ;
  513 :out<= 0 ;
  514 :out<= 0 ;
  515 :out<= 0 ;
  516 :out<= 0 ;
  517 :out<= 0 ;
  518 :out<= 0 ;
  519 :out<= 0 ;
  520 :out<= 0 ;
  521 :out<= 0 ;
  522 :out<= 0 ;
  523 :out<= 0 ;
  524 :out<= 0 ;
  525 :out<= 0 ;
  526 :out<= 0 ;
  527 :out<= 0 ;
  528 :out<= 0 ;
  529 :out<= 0 ;
  530 :out<= 0 ;
  531 :out<= 0 ;
  532 :out<= 0 ;
  533 :out<= 0 ;
  534 :out<= 0 ;
  535 :out<= 0 ;
  536 :out<= 0 ;
  537 :out<= 0 ;
  538 :out<= 0 ;
  539 :out<= 0 ;
  540 :out<= 0 ;
  541 :out<= 0 ;
  542 :out<= 0 ;
  543 :out<= 0 ;
  544 :out<= 0 ;
  545 :out<= 0 ;
  546 :out<= 0 ;
  547 :out<= 0 ;
  548 :out<= 0 ;
  549 :out<= 0 ;
  550 :out<= 0 ;
  551 :out<= 0 ;
  552 :out<= 0 ;
  553 :out<= 0 ;
  554 :out<= 0 ;
  555 :out<= 0 ;
  556 :out<= 0 ;
  557 :out<= 0 ;
  558 :out<= 0 ;
  559 :out<= 1 ;
  560 :out<= 0 ;
  561 :out<= 0 ;
  562 :out<= 0 ;
  563 :out<= 0 ;
  564 :out<= 0 ;
  565 :out<= 0 ;
  566 :out<= 0 ;
  567 :out<= 1 ;
  568 :out<= 0 ;
  569 :out<= 0 ;
  570 :out<= 0 ;
  571 :out<= 1 ;
  572 :out<= 0 ;
  573 :out<= 1 ;
  574 :out<= 1 ;
  575 :out<= 1 ;
  576 :out<= 0 ;
  577 :out<= 0 ;
  578 :out<= 0 ;
  579 :out<= 0 ;
  580 :out<= 0 ;
  581 :out<= 0 ;
  582 :out<= 0 ;
  583 :out<= 0 ;
  584 :out<= 0 ;
  585 :out<= 0 ;
  586 :out<= 0 ;
  587 :out<= 0 ;
  588 :out<= 0 ;
  589 :out<= 0 ;
  590 :out<= 0 ;
  591 :out<= 1 ;
  592 :out<= 0 ;
  593 :out<= 0 ;
  594 :out<= 0 ;
  595 :out<= 0 ;
  596 :out<= 0 ;
  597 :out<= 1 ;
  598 :out<= 1 ;
  599 :out<= 1 ;
  600 :out<= 0 ;
  601 :out<= 1 ;
  602 :out<= 1 ;
  603 :out<= 1 ;
  604 :out<= 1 ;
  605 :out<= 1 ;
  606 :out<= 1 ;
  607 :out<= 1 ;
  608 :out<= 0 ;
  609 :out<= 0 ;
  610 :out<= 0 ;
  611 :out<= 1 ;
  612 :out<= 0 ;
  613 :out<= 1 ;
  614 :out<= 1 ;
  615 :out<= 1 ;
  616 :out<= 0 ;
  617 :out<= 1 ;
  618 :out<= 1 ;
  619 :out<= 1 ;
  620 :out<= 1 ;
  621 :out<= 1 ;
  622 :out<= 1 ;
  623 :out<= 1 ;
  624 :out<= 0 ;
  625 :out<= 1 ;
  626 :out<= 1 ;
  627 :out<= 1 ;
  628 :out<= 1 ;
  629 :out<= 1 ;
  630 :out<= 1 ;
  631 :out<= 1 ;
  632 :out<= 1 ;
  633 :out<= 1 ;
  634 :out<= 1 ;
  635 :out<= 1 ;
  636 :out<= 1 ;
  637 :out<= 1 ;
  638 :out<= 1 ;
  639 :out<= 1 ;
  640 :out<= 0 ;
  641 :out<= 0 ;
  642 :out<= 0 ;
  643 :out<= 0 ;
  644 :out<= 0 ;
  645 :out<= 0 ;
  646 :out<= 0 ;
  647 :out<= 0 ;
  648 :out<= 0 ;
  649 :out<= 0 ;
  650 :out<= 0 ;
  651 :out<= 1 ;
  652 :out<= 0 ;
  653 :out<= 1 ;
  654 :out<= 1 ;
  655 :out<= 1 ;
  656 :out<= 0 ;
  657 :out<= 0 ;
  658 :out<= 0 ;
  659 :out<= 1 ;
  660 :out<= 0 ;
  661 :out<= 1 ;
  662 :out<= 1 ;
  663 :out<= 1 ;
  664 :out<= 0 ;
  665 :out<= 1 ;
  666 :out<= 1 ;
  667 :out<= 1 ;
  668 :out<= 1 ;
  669 :out<= 1 ;
  670 :out<= 1 ;
  671 :out<= 1 ;
  672 :out<= 0 ;
  673 :out<= 0 ;
  674 :out<= 0 ;
  675 :out<= 1 ;
  676 :out<= 0 ;
  677 :out<= 1 ;
  678 :out<= 1 ;
  679 :out<= 1 ;
  680 :out<= 0 ;
  681 :out<= 1 ;
  682 :out<= 1 ;
  683 :out<= 1 ;
  684 :out<= 1 ;
  685 :out<= 1 ;
  686 :out<= 1 ;
  687 :out<= 1 ;
  688 :out<= 0 ;
  689 :out<= 1 ;
  690 :out<= 1 ;
  691 :out<= 1 ;
  692 :out<= 1 ;
  693 :out<= 1 ;
  694 :out<= 1 ;
  695 :out<= 1 ;
  696 :out<= 1 ;
  697 :out<= 1 ;
  698 :out<= 1 ;
  699 :out<= 1 ;
  700 :out<= 1 ;
  701 :out<= 1 ;
  702 :out<= 1 ;
  703 :out<= 1 ;
  704 :out<= 0 ;
  705 :out<= 0 ;
  706 :out<= 0 ;
  707 :out<= 1 ;
  708 :out<= 0 ;
  709 :out<= 1 ;
  710 :out<= 1 ;
  711 :out<= 1 ;
  712 :out<= 0 ;
  713 :out<= 1 ;
  714 :out<= 1 ;
  715 :out<= 1 ;
  716 :out<= 1 ;
  717 :out<= 1 ;
  718 :out<= 1 ;
  719 :out<= 1 ;
  720 :out<= 1 ;
  721 :out<= 1 ;
  722 :out<= 1 ;
  723 :out<= 1 ;
  724 :out<= 1 ;
  725 :out<= 1 ;
  726 :out<= 1 ;
  727 :out<= 1 ;
  728 :out<= 1 ;
  729 :out<= 1 ;
  730 :out<= 1 ;
  731 :out<= 1 ;
  732 :out<= 1 ;
  733 :out<= 1 ;
  734 :out<= 1 ;
  735 :out<= 1 ;
  736 :out<= 1 ;
  737 :out<= 1 ;
  738 :out<= 1 ;
  739 :out<= 1 ;
  740 :out<= 1 ;
  741 :out<= 1 ;
  742 :out<= 1 ;
  743 :out<= 1 ;
  744 :out<= 1 ;
  745 :out<= 1 ;
  746 :out<= 1 ;
  747 :out<= 1 ;
  748 :out<= 1 ;
  749 :out<= 1 ;
  750 :out<= 1 ;
  751 :out<= 1 ;
  752 :out<= 1 ;
  753 :out<= 1 ;
  754 :out<= 1 ;
  755 :out<= 1 ;
  756 :out<= 1 ;
  757 :out<= 1 ;
  758 :out<= 1 ;
  759 :out<= 1 ;
  760 :out<= 1 ;
  761 :out<= 1 ;
  762 :out<= 1 ;
  763 :out<= 1 ;
  764 :out<= 1 ;
  765 :out<= 1 ;
  766 :out<= 1 ;
  767 :out<= 1 ;
  768 :out<= 0 ;
  769 :out<= 0 ;
  770 :out<= 0 ;
  771 :out<= 0 ;
  772 :out<= 0 ;
  773 :out<= 0 ;
  774 :out<= 0 ;
  775 :out<= 1 ;
  776 :out<= 0 ;
  777 :out<= 0 ;
  778 :out<= 0 ;
  779 :out<= 1 ;
  780 :out<= 0 ;
  781 :out<= 1 ;
  782 :out<= 1 ;
  783 :out<= 1 ;
  784 :out<= 0 ;
  785 :out<= 0 ;
  786 :out<= 0 ;
  787 :out<= 1 ;
  788 :out<= 0 ;
  789 :out<= 1 ;
  790 :out<= 1 ;
  791 :out<= 1 ;
  792 :out<= 0 ;
  793 :out<= 1 ;
  794 :out<= 1 ;
  795 :out<= 1 ;
  796 :out<= 1 ;
  797 :out<= 1 ;
  798 :out<= 1 ;
  799 :out<= 1 ;
  800 :out<= 0 ;
  801 :out<= 0 ;
  802 :out<= 0 ;
  803 :out<= 1 ;
  804 :out<= 1 ;
  805 :out<= 1 ;
  806 :out<= 1 ;
  807 :out<= 1 ;
  808 :out<= 1 ;
  809 :out<= 1 ;
  810 :out<= 1 ;
  811 :out<= 1 ;
  812 :out<= 1 ;
  813 :out<= 1 ;
  814 :out<= 1 ;
  815 :out<= 1 ;
  816 :out<= 1 ;
  817 :out<= 1 ;
  818 :out<= 1 ;
  819 :out<= 1 ;
  820 :out<= 1 ;
  821 :out<= 1 ;
  822 :out<= 1 ;
  823 :out<= 1 ;
  824 :out<= 1 ;
  825 :out<= 1 ;
  826 :out<= 1 ;
  827 :out<= 1 ;
  828 :out<= 1 ;
  829 :out<= 1 ;
  830 :out<= 1 ;
  831 :out<= 1 ;
  832 :out<= 0 ;
  833 :out<= 0 ;
  834 :out<= 1 ;
  835 :out<= 1 ;
  836 :out<= 1 ;
  837 :out<= 1 ;
  838 :out<= 1 ;
  839 :out<= 1 ;
  840 :out<= 1 ;
  841 :out<= 1 ;
  842 :out<= 1 ;
  843 :out<= 1 ;
  844 :out<= 1 ;
  845 :out<= 1 ;
  846 :out<= 1 ;
  847 :out<= 1 ;
  848 :out<= 1 ;
  849 :out<= 1 ;
  850 :out<= 1 ;
  851 :out<= 1 ;
  852 :out<= 1 ;
  853 :out<= 1 ;
  854 :out<= 1 ;
  855 :out<= 1 ;
  856 :out<= 1 ;
  857 :out<= 1 ;
  858 :out<= 1 ;
  859 :out<= 1 ;
  860 :out<= 1 ;
  861 :out<= 1 ;
  862 :out<= 1 ;
  863 :out<= 1 ;
  864 :out<= 1 ;
  865 :out<= 1 ;
  866 :out<= 1 ;
  867 :out<= 1 ;
  868 :out<= 1 ;
  869 :out<= 1 ;
  870 :out<= 1 ;
  871 :out<= 1 ;
  872 :out<= 1 ;
  873 :out<= 1 ;
  874 :out<= 1 ;
  875 :out<= 1 ;
  876 :out<= 1 ;
  877 :out<= 1 ;
  878 :out<= 1 ;
  879 :out<= 1 ;
  880 :out<= 1 ;
  881 :out<= 1 ;
  882 :out<= 1 ;
  883 :out<= 1 ;
  884 :out<= 1 ;
  885 :out<= 1 ;
  886 :out<= 1 ;
  887 :out<= 1 ;
  888 :out<= 1 ;
  889 :out<= 1 ;
  890 :out<= 1 ;
  891 :out<= 1 ;
  892 :out<= 1 ;
  893 :out<= 1 ;
  894 :out<= 1 ;
  895 :out<= 1 ;
  896 :out<= 0 ;
  897 :out<= 1 ;
  898 :out<= 1 ;
  899 :out<= 1 ;
  900 :out<= 1 ;
  901 :out<= 1 ;
  902 :out<= 1 ;
  903 :out<= 1 ;
  904 :out<= 1 ;
  905 :out<= 1 ;
  906 :out<= 1 ;
  907 :out<= 1 ;
  908 :out<= 1 ;
  909 :out<= 1 ;
  910 :out<= 1 ;
  911 :out<= 1 ;
  912 :out<= 1 ;
  913 :out<= 1 ;
  914 :out<= 1 ;
  915 :out<= 1 ;
  916 :out<= 1 ;
  917 :out<= 1 ;
  918 :out<= 1 ;
  919 :out<= 1 ;
  920 :out<= 1 ;
  921 :out<= 1 ;
  922 :out<= 1 ;
  923 :out<= 1 ;
  924 :out<= 1 ;
  925 :out<= 1 ;
  926 :out<= 1 ;
  927 :out<= 1 ;
  928 :out<= 1 ;
  929 :out<= 1 ;
  930 :out<= 1 ;
  931 :out<= 1 ;
  932 :out<= 1 ;
  933 :out<= 1 ;
  934 :out<= 1 ;
  935 :out<= 1 ;
  936 :out<= 1 ;
  937 :out<= 1 ;
  938 :out<= 1 ;
  939 :out<= 1 ;
  940 :out<= 1 ;
  941 :out<= 1 ;
  942 :out<= 1 ;
  943 :out<= 1 ;
  944 :out<= 1 ;
  945 :out<= 1 ;
  946 :out<= 1 ;
  947 :out<= 1 ;
  948 :out<= 1 ;
  949 :out<= 1 ;
  950 :out<= 1 ;
  951 :out<= 1 ;
  952 :out<= 1 ;
  953 :out<= 1 ;
  954 :out<= 1 ;
  955 :out<= 1 ;
  956 :out<= 1 ;
  957 :out<= 1 ;
  958 :out<= 1 ;
  959 :out<= 1 ;
  960 :out<= 1 ;
  961 :out<= 1 ;
  962 :out<= 1 ;
  963 :out<= 1 ;
  964 :out<= 1 ;
  965 :out<= 1 ;
  966 :out<= 1 ;
  967 :out<= 1 ;
  968 :out<= 1 ;
  969 :out<= 1 ;
  970 :out<= 1 ;
  971 :out<= 1 ;
  972 :out<= 1 ;
  973 :out<= 1 ;
  974 :out<= 1 ;
  975 :out<= 1 ;
  976 :out<= 1 ;
  977 :out<= 1 ;
  978 :out<= 1 ;
  979 :out<= 1 ;
  980 :out<= 1 ;
  981 :out<= 1 ;
  982 :out<= 1 ;
  983 :out<= 1 ;
  984 :out<= 1 ;
  985 :out<= 1 ;
  986 :out<= 1 ;
  987 :out<= 1 ;
  988 :out<= 1 ;
  989 :out<= 1 ;
  990 :out<= 1 ;
  991 :out<= 1 ;
  992 :out<= 1 ;
  993 :out<= 1 ;
  994 :out<= 1 ;
  995 :out<= 1 ;
  996 :out<= 1 ;
  997 :out<= 1 ;
  998 :out<= 1 ;
  999 :out<= 1 ;
  1000 :out<= 1 ;
  1001 :out<= 1 ;
  1002 :out<= 1 ;
  1003 :out<= 1 ;
  1004 :out<= 1 ;
  1005 :out<= 1 ;
  1006 :out<= 1 ;
  1007 :out<= 1 ;
  1008 :out<= 1 ;
  1009 :out<= 1 ;
  1010 :out<= 1 ;
  1011 :out<= 1 ;
  1012 :out<= 1 ;
  1013 :out<= 1 ;
  1014 :out<= 1 ;
  1015 :out<= 1 ;
  1016 :out<= 1 ;
  1017 :out<= 1 ;
  1018 :out<= 1 ;
  1019 :out<= 1 ;
  1020 :out<= 1 ;
  1021 :out<= 1 ;
  1022 :out<= 1 ;
  1023 :out<= 1 ;
 endcase
case(in_bit_index2)
  0 :out2<= 0 ;
  1 :out2<= 0 ;
  2 :out2<= 0 ;
  3 :out2<= 0 ;
  4 :out2<= 0 ;
  5 :out2<= 0 ;
  6 :out2<= 0 ;
  7 :out2<= 0 ;
  8 :out2<= 0 ;
  9 :out2<= 0 ;
  10 :out2<= 0 ;
  11 :out2<= 0 ;
  12 :out2<= 0 ;
  13 :out2<= 0 ;
  14 :out2<= 0 ;
  15 :out2<= 0 ;
  16 :out2<= 0 ;
  17 :out2<= 0 ;
  18 :out2<= 0 ;
  19 :out2<= 0 ;
  20 :out2<= 0 ;
  21 :out2<= 0 ;
  22 :out2<= 0 ;
  23 :out2<= 0 ;
  24 :out2<= 0 ;
  25 :out2<= 0 ;
  26 :out2<= 0 ;
  27 :out2<= 0 ;
  28 :out2<= 0 ;
  29 :out2<= 0 ;
  30 :out2<= 0 ;
  31 :out2<= 0 ;
  32 :out2<= 0 ;
  33 :out2<= 0 ;
  34 :out2<= 0 ;
  35 :out2<= 0 ;
  36 :out2<= 0 ;
  37 :out2<= 0 ;
  38 :out2<= 0 ;
  39 :out2<= 0 ;
  40 :out2<= 0 ;
  41 :out2<= 0 ;
  42 :out2<= 0 ;
  43 :out2<= 0 ;
  44 :out2<= 0 ;
  45 :out2<= 0 ;
  46 :out2<= 0 ;
  47 :out2<= 0 ;
  48 :out2<= 0 ;
  49 :out2<= 0 ;
  50 :out2<= 0 ;
  51 :out2<= 0 ;
  52 :out2<= 0 ;
  53 :out2<= 0 ;
  54 :out2<= 0 ;
  55 :out2<= 0 ;
  56 :out2<= 0 ;
  57 :out2<= 0 ;
  58 :out2<= 0 ;
  59 :out2<= 0 ;
  60 :out2<= 0 ;
  61 :out2<= 0 ;
  62 :out2<= 0 ;
  63 :out2<= 0 ;
  64 :out2<= 0 ;
  65 :out2<= 0 ;
  66 :out2<= 0 ;
  67 :out2<= 0 ;
  68 :out2<= 0 ;
  69 :out2<= 0 ;
  70 :out2<= 0 ;
  71 :out2<= 0 ;
  72 :out2<= 0 ;
  73 :out2<= 0 ;
  74 :out2<= 0 ;
  75 :out2<= 0 ;
  76 :out2<= 0 ;
  77 :out2<= 0 ;
  78 :out2<= 0 ;
  79 :out2<= 0 ;
  80 :out2<= 0 ;
  81 :out2<= 0 ;
  82 :out2<= 0 ;
  83 :out2<= 0 ;
  84 :out2<= 0 ;
  85 :out2<= 0 ;
  86 :out2<= 0 ;
  87 :out2<= 0 ;
  88 :out2<= 0 ;
  89 :out2<= 0 ;
  90 :out2<= 0 ;
  91 :out2<= 0 ;
  92 :out2<= 0 ;
  93 :out2<= 0 ;
  94 :out2<= 0 ;
  95 :out2<= 0 ;
  96 :out2<= 0 ;
  97 :out2<= 0 ;
  98 :out2<= 0 ;
  99 :out2<= 0 ;
  100 :out2<= 0 ;
  101 :out2<= 0 ;
  102 :out2<= 0 ;
  103 :out2<= 0 ;
  104 :out2<= 0 ;
  105 :out2<= 0 ;
  106 :out2<= 0 ;
  107 :out2<= 0 ;
  108 :out2<= 0 ;
  109 :out2<= 0 ;
  110 :out2<= 0 ;
  111 :out2<= 0 ;
  112 :out2<= 0 ;
  113 :out2<= 0 ;
  114 :out2<= 0 ;
  115 :out2<= 0 ;
  116 :out2<= 0 ;
  117 :out2<= 0 ;
  118 :out2<= 0 ;
  119 :out2<= 0 ;
  120 :out2<= 0 ;
  121 :out2<= 0 ;
  122 :out2<= 0 ;
  123 :out2<= 0 ;
  124 :out2<= 0 ;
  125 :out2<= 0 ;
  126 :out2<= 0 ;
  127 :out2<= 0 ;
  128 :out2<= 0 ;
  129 :out2<= 0 ;
  130 :out2<= 0 ;
  131 :out2<= 0 ;
  132 :out2<= 0 ;
  133 :out2<= 0 ;
  134 :out2<= 0 ;
  135 :out2<= 0 ;
  136 :out2<= 0 ;
  137 :out2<= 0 ;
  138 :out2<= 0 ;
  139 :out2<= 0 ;
  140 :out2<= 0 ;
  141 :out2<= 0 ;
  142 :out2<= 0 ;
  143 :out2<= 0 ;
  144 :out2<= 0 ;
  145 :out2<= 0 ;
  146 :out2<= 0 ;
  147 :out2<= 0 ;
  148 :out2<= 0 ;
  149 :out2<= 0 ;
  150 :out2<= 0 ;
  151 :out2<= 0 ;
  152 :out2<= 0 ;
  153 :out2<= 0 ;
  154 :out2<= 0 ;
  155 :out2<= 0 ;
  156 :out2<= 0 ;
  157 :out2<= 0 ;
  158 :out2<= 0 ;
  159 :out2<= 0 ;
  160 :out2<= 0 ;
  161 :out2<= 0 ;
  162 :out2<= 0 ;
  163 :out2<= 0 ;
  164 :out2<= 0 ;
  165 :out2<= 0 ;
  166 :out2<= 0 ;
  167 :out2<= 0 ;
  168 :out2<= 0 ;
  169 :out2<= 0 ;
  170 :out2<= 0 ;
  171 :out2<= 0 ;
  172 :out2<= 0 ;
  173 :out2<= 0 ;
  174 :out2<= 0 ;
  175 :out2<= 0 ;
  176 :out2<= 0 ;
  177 :out2<= 0 ;
  178 :out2<= 0 ;
  179 :out2<= 0 ;
  180 :out2<= 0 ;
  181 :out2<= 0 ;
  182 :out2<= 0 ;
  183 :out2<= 0 ;
  184 :out2<= 0 ;
  185 :out2<= 0 ;
  186 :out2<= 0 ;
  187 :out2<= 0 ;
  188 :out2<= 0 ;
  189 :out2<= 0 ;
  190 :out2<= 0 ;
  191 :out2<= 1 ;
  192 :out2<= 0 ;
  193 :out2<= 0 ;
  194 :out2<= 0 ;
  195 :out2<= 0 ;
  196 :out2<= 0 ;
  197 :out2<= 0 ;
  198 :out2<= 0 ;
  199 :out2<= 0 ;
  200 :out2<= 0 ;
  201 :out2<= 0 ;
  202 :out2<= 0 ;
  203 :out2<= 0 ;
  204 :out2<= 0 ;
  205 :out2<= 0 ;
  206 :out2<= 0 ;
  207 :out2<= 0 ;
  208 :out2<= 0 ;
  209 :out2<= 0 ;
  210 :out2<= 0 ;
  211 :out2<= 0 ;
  212 :out2<= 0 ;
  213 :out2<= 0 ;
  214 :out2<= 0 ;
  215 :out2<= 0 ;
  216 :out2<= 0 ;
  217 :out2<= 0 ;
  218 :out2<= 0 ;
  219 :out2<= 0 ;
  220 :out2<= 0 ;
  221 :out2<= 0 ;
  222 :out2<= 0 ;
  223 :out2<= 1 ;
  224 :out2<= 0 ;
  225 :out2<= 0 ;
  226 :out2<= 0 ;
  227 :out2<= 0 ;
  228 :out2<= 0 ;
  229 :out2<= 0 ;
  230 :out2<= 0 ;
  231 :out2<= 0 ;
  232 :out2<= 0 ;
  233 :out2<= 0 ;
  234 :out2<= 0 ;
  235 :out2<= 1 ;
  236 :out2<= 0 ;
  237 :out2<= 1 ;
  238 :out2<= 1 ;
  239 :out2<= 1 ;
  240 :out2<= 0 ;
  241 :out2<= 0 ;
  242 :out2<= 0 ;
  243 :out2<= 1 ;
  244 :out2<= 0 ;
  245 :out2<= 1 ;
  246 :out2<= 1 ;
  247 :out2<= 1 ;
  248 :out2<= 0 ;
  249 :out2<= 1 ;
  250 :out2<= 1 ;
  251 :out2<= 1 ;
  252 :out2<= 1 ;
  253 :out2<= 1 ;
  254 :out2<= 1 ;
  255 :out2<= 1 ;
  256 :out2<= 0 ;
  257 :out2<= 0 ;
  258 :out2<= 0 ;
  259 :out2<= 0 ;
  260 :out2<= 0 ;
  261 :out2<= 0 ;
  262 :out2<= 0 ;
  263 :out2<= 0 ;
  264 :out2<= 0 ;
  265 :out2<= 0 ;
  266 :out2<= 0 ;
  267 :out2<= 0 ;
  268 :out2<= 0 ;
  269 :out2<= 0 ;
  270 :out2<= 0 ;
  271 :out2<= 0 ;
  272 :out2<= 0 ;
  273 :out2<= 0 ;
  274 :out2<= 0 ;
  275 :out2<= 0 ;
  276 :out2<= 0 ;
  277 :out2<= 0 ;
  278 :out2<= 0 ;
  279 :out2<= 0 ;
  280 :out2<= 0 ;
  281 :out2<= 0 ;
  282 :out2<= 0 ;
  283 :out2<= 0 ;
  284 :out2<= 0 ;
  285 :out2<= 0 ;
  286 :out2<= 0 ;
  287 :out2<= 0 ;
  288 :out2<= 0 ;
  289 :out2<= 0 ;
  290 :out2<= 0 ;
  291 :out2<= 0 ;
  292 :out2<= 0 ;
  293 :out2<= 0 ;
  294 :out2<= 0 ;
  295 :out2<= 0 ;
  296 :out2<= 0 ;
  297 :out2<= 0 ;
  298 :out2<= 0 ;
  299 :out2<= 0 ;
  300 :out2<= 0 ;
  301 :out2<= 0 ;
  302 :out2<= 0 ;
  303 :out2<= 0 ;
  304 :out2<= 0 ;
  305 :out2<= 0 ;
  306 :out2<= 0 ;
  307 :out2<= 0 ;
  308 :out2<= 0 ;
  309 :out2<= 0 ;
  310 :out2<= 0 ;
  311 :out2<= 0 ;
  312 :out2<= 0 ;
  313 :out2<= 0 ;
  314 :out2<= 0 ;
  315 :out2<= 1 ;
  316 :out2<= 0 ;
  317 :out2<= 1 ;
  318 :out2<= 1 ;
  319 :out2<= 1 ;
  320 :out2<= 0 ;
  321 :out2<= 0 ;
  322 :out2<= 0 ;
  323 :out2<= 0 ;
  324 :out2<= 0 ;
  325 :out2<= 0 ;
  326 :out2<= 0 ;
  327 :out2<= 0 ;
  328 :out2<= 0 ;
  329 :out2<= 0 ;
  330 :out2<= 0 ;
  331 :out2<= 0 ;
  332 :out2<= 0 ;
  333 :out2<= 0 ;
  334 :out2<= 0 ;
  335 :out2<= 0 ;
  336 :out2<= 0 ;
  337 :out2<= 0 ;
  338 :out2<= 0 ;
  339 :out2<= 0 ;
  340 :out2<= 0 ;
  341 :out2<= 0 ;
  342 :out2<= 0 ;
  343 :out2<= 1 ;
  344 :out2<= 0 ;
  345 :out2<= 0 ;
  346 :out2<= 0 ;
  347 :out2<= 1 ;
  348 :out2<= 0 ;
  349 :out2<= 1 ;
  350 :out2<= 1 ;
  351 :out2<= 1 ;
  352 :out2<= 0 ;
  353 :out2<= 0 ;
  354 :out2<= 0 ;
  355 :out2<= 0 ;
  356 :out2<= 0 ;
  357 :out2<= 0 ;
  358 :out2<= 0 ;
  359 :out2<= 1 ;
  360 :out2<= 0 ;
  361 :out2<= 0 ;
  362 :out2<= 0 ;
  363 :out2<= 1 ;
  364 :out2<= 0 ;
  365 :out2<= 1 ;
  366 :out2<= 1 ;
  367 :out2<= 1 ;
  368 :out2<= 0 ;
  369 :out2<= 0 ;
  370 :out2<= 1 ;
  371 :out2<= 1 ;
  372 :out2<= 1 ;
  373 :out2<= 1 ;
  374 :out2<= 1 ;
  375 :out2<= 1 ;
  376 :out2<= 1 ;
  377 :out2<= 1 ;
  378 :out2<= 1 ;
  379 :out2<= 1 ;
  380 :out2<= 1 ;
  381 :out2<= 1 ;
  382 :out2<= 1 ;
  383 :out2<= 1 ;
  384 :out2<= 0 ;
  385 :out2<= 0 ;
  386 :out2<= 0 ;
  387 :out2<= 0 ;
  388 :out2<= 0 ;
  389 :out2<= 0 ;
  390 :out2<= 0 ;
  391 :out2<= 0 ;
  392 :out2<= 0 ;
  393 :out2<= 0 ;
  394 :out2<= 0 ;
  395 :out2<= 0 ;
  396 :out2<= 0 ;
  397 :out2<= 0 ;
  398 :out2<= 0 ;
  399 :out2<= 1 ;
  400 :out2<= 0 ;
  401 :out2<= 0 ;
  402 :out2<= 0 ;
  403 :out2<= 0 ;
  404 :out2<= 0 ;
  405 :out2<= 0 ;
  406 :out2<= 0 ;
  407 :out2<= 1 ;
  408 :out2<= 0 ;
  409 :out2<= 0 ;
  410 :out2<= 1 ;
  411 :out2<= 1 ;
  412 :out2<= 1 ;
  413 :out2<= 1 ;
  414 :out2<= 1 ;
  415 :out2<= 1 ;
  416 :out2<= 0 ;
  417 :out2<= 0 ;
  418 :out2<= 0 ;
  419 :out2<= 0 ;
  420 :out2<= 0 ;
  421 :out2<= 1 ;
  422 :out2<= 1 ;
  423 :out2<= 1 ;
  424 :out2<= 0 ;
  425 :out2<= 1 ;
  426 :out2<= 1 ;
  427 :out2<= 1 ;
  428 :out2<= 1 ;
  429 :out2<= 1 ;
  430 :out2<= 1 ;
  431 :out2<= 1 ;
  432 :out2<= 0 ;
  433 :out2<= 1 ;
  434 :out2<= 1 ;
  435 :out2<= 1 ;
  436 :out2<= 1 ;
  437 :out2<= 1 ;
  438 :out2<= 1 ;
  439 :out2<= 1 ;
  440 :out2<= 1 ;
  441 :out2<= 1 ;
  442 :out2<= 1 ;
  443 :out2<= 1 ;
  444 :out2<= 1 ;
  445 :out2<= 1 ;
  446 :out2<= 1 ;
  447 :out2<= 1 ;
  448 :out2<= 0 ;
  449 :out2<= 0 ;
  450 :out2<= 0 ;
  451 :out2<= 1 ;
  452 :out2<= 0 ;
  453 :out2<= 1 ;
  454 :out2<= 1 ;
  455 :out2<= 1 ;
  456 :out2<= 0 ;
  457 :out2<= 1 ;
  458 :out2<= 1 ;
  459 :out2<= 1 ;
  460 :out2<= 1 ;
  461 :out2<= 1 ;
  462 :out2<= 1 ;
  463 :out2<= 1 ;
  464 :out2<= 0 ;
  465 :out2<= 1 ;
  466 :out2<= 1 ;
  467 :out2<= 1 ;
  468 :out2<= 1 ;
  469 :out2<= 1 ;
  470 :out2<= 1 ;
  471 :out2<= 1 ;
  472 :out2<= 1 ;
  473 :out2<= 1 ;
  474 :out2<= 1 ;
  475 :out2<= 1 ;
  476 :out2<= 1 ;
  477 :out2<= 1 ;
  478 :out2<= 1 ;
  479 :out2<= 1 ;
  480 :out2<= 0 ;
  481 :out2<= 1 ;
  482 :out2<= 1 ;
  483 :out2<= 1 ;
  484 :out2<= 1 ;
  485 :out2<= 1 ;
  486 :out2<= 1 ;
  487 :out2<= 1 ;
  488 :out2<= 1 ;
  489 :out2<= 1 ;
  490 :out2<= 1 ;
  491 :out2<= 1 ;
  492 :out2<= 1 ;
  493 :out2<= 1 ;
  494 :out2<= 1 ;
  495 :out2<= 1 ;
  496 :out2<= 1 ;
  497 :out2<= 1 ;
  498 :out2<= 1 ;
  499 :out2<= 1 ;
  500 :out2<= 1 ;
  501 :out2<= 1 ;
  502 :out2<= 1 ;
  503 :out2<= 1 ;
  504 :out2<= 1 ;
  505 :out2<= 1 ;
  506 :out2<= 1 ;
  507 :out2<= 1 ;
  508 :out2<= 1 ;
  509 :out2<= 1 ;
  510 :out2<= 1 ;
  511 :out2<= 1 ;
  512 :out2<= 0 ;
  513 :out2<= 0 ;
  514 :out2<= 0 ;
  515 :out2<= 0 ;
  516 :out2<= 0 ;
  517 :out2<= 0 ;
  518 :out2<= 0 ;
  519 :out2<= 0 ;
  520 :out2<= 0 ;
  521 :out2<= 0 ;
  522 :out2<= 0 ;
  523 :out2<= 0 ;
  524 :out2<= 0 ;
  525 :out2<= 0 ;
  526 :out2<= 0 ;
  527 :out2<= 0 ;
  528 :out2<= 0 ;
  529 :out2<= 0 ;
  530 :out2<= 0 ;
  531 :out2<= 0 ;
  532 :out2<= 0 ;
  533 :out2<= 0 ;
  534 :out2<= 0 ;
  535 :out2<= 0 ;
  536 :out2<= 0 ;
  537 :out2<= 0 ;
  538 :out2<= 0 ;
  539 :out2<= 0 ;
  540 :out2<= 0 ;
  541 :out2<= 0 ;
  542 :out2<= 0 ;
  543 :out2<= 0 ;
  544 :out2<= 0 ;
  545 :out2<= 0 ;
  546 :out2<= 0 ;
  547 :out2<= 0 ;
  548 :out2<= 0 ;
  549 :out2<= 0 ;
  550 :out2<= 0 ;
  551 :out2<= 0 ;
  552 :out2<= 0 ;
  553 :out2<= 0 ;
  554 :out2<= 0 ;
  555 :out2<= 0 ;
  556 :out2<= 0 ;
  557 :out2<= 0 ;
  558 :out2<= 0 ;
  559 :out2<= 1 ;
  560 :out2<= 0 ;
  561 :out2<= 0 ;
  562 :out2<= 0 ;
  563 :out2<= 0 ;
  564 :out2<= 0 ;
  565 :out2<= 0 ;
  566 :out2<= 0 ;
  567 :out2<= 1 ;
  568 :out2<= 0 ;
  569 :out2<= 0 ;
  570 :out2<= 0 ;
  571 :out2<= 1 ;
  572 :out2<= 0 ;
  573 :out2<= 1 ;
  574 :out2<= 1 ;
  575 :out2<= 1 ;
  576 :out2<= 0 ;
  577 :out2<= 0 ;
  578 :out2<= 0 ;
  579 :out2<= 0 ;
  580 :out2<= 0 ;
  581 :out2<= 0 ;
  582 :out2<= 0 ;
  583 :out2<= 0 ;
  584 :out2<= 0 ;
  585 :out2<= 0 ;
  586 :out2<= 0 ;
  587 :out2<= 0 ;
  588 :out2<= 0 ;
  589 :out2<= 0 ;
  590 :out2<= 0 ;
  591 :out2<= 1 ;
  592 :out2<= 0 ;
  593 :out2<= 0 ;
  594 :out2<= 0 ;
  595 :out2<= 0 ;
  596 :out2<= 0 ;
  597 :out2<= 1 ;
  598 :out2<= 1 ;
  599 :out2<= 1 ;
  600 :out2<= 0 ;
  601 :out2<= 1 ;
  602 :out2<= 1 ;
  603 :out2<= 1 ;
  604 :out2<= 1 ;
  605 :out2<= 1 ;
  606 :out2<= 1 ;
  607 :out2<= 1 ;
  608 :out2<= 0 ;
  609 :out2<= 0 ;
  610 :out2<= 0 ;
  611 :out2<= 1 ;
  612 :out2<= 0 ;
  613 :out2<= 1 ;
  614 :out2<= 1 ;
  615 :out2<= 1 ;
  616 :out2<= 0 ;
  617 :out2<= 1 ;
  618 :out2<= 1 ;
  619 :out2<= 1 ;
  620 :out2<= 1 ;
  621 :out2<= 1 ;
  622 :out2<= 1 ;
  623 :out2<= 1 ;
  624 :out2<= 0 ;
  625 :out2<= 1 ;
  626 :out2<= 1 ;
  627 :out2<= 1 ;
  628 :out2<= 1 ;
  629 :out2<= 1 ;
  630 :out2<= 1 ;
  631 :out2<= 1 ;
  632 :out2<= 1 ;
  633 :out2<= 1 ;
  634 :out2<= 1 ;
  635 :out2<= 1 ;
  636 :out2<= 1 ;
  637 :out2<= 1 ;
  638 :out2<= 1 ;
  639 :out2<= 1 ;
  640 :out2<= 0 ;
  641 :out2<= 0 ;
  642 :out2<= 0 ;
  643 :out2<= 0 ;
  644 :out2<= 0 ;
  645 :out2<= 0 ;
  646 :out2<= 0 ;
  647 :out2<= 0 ;
  648 :out2<= 0 ;
  649 :out2<= 0 ;
  650 :out2<= 0 ;
  651 :out2<= 1 ;
  652 :out2<= 0 ;
  653 :out2<= 1 ;
  654 :out2<= 1 ;
  655 :out2<= 1 ;
  656 :out2<= 0 ;
  657 :out2<= 0 ;
  658 :out2<= 0 ;
  659 :out2<= 1 ;
  660 :out2<= 0 ;
  661 :out2<= 1 ;
  662 :out2<= 1 ;
  663 :out2<= 1 ;
  664 :out2<= 0 ;
  665 :out2<= 1 ;
  666 :out2<= 1 ;
  667 :out2<= 1 ;
  668 :out2<= 1 ;
  669 :out2<= 1 ;
  670 :out2<= 1 ;
  671 :out2<= 1 ;
  672 :out2<= 0 ;
  673 :out2<= 0 ;
  674 :out2<= 0 ;
  675 :out2<= 1 ;
  676 :out2<= 0 ;
  677 :out2<= 1 ;
  678 :out2<= 1 ;
  679 :out2<= 1 ;
  680 :out2<= 0 ;
  681 :out2<= 1 ;
  682 :out2<= 1 ;
  683 :out2<= 1 ;
  684 :out2<= 1 ;
  685 :out2<= 1 ;
  686 :out2<= 1 ;
  687 :out2<= 1 ;
  688 :out2<= 0 ;
  689 :out2<= 1 ;
  690 :out2<= 1 ;
  691 :out2<= 1 ;
  692 :out2<= 1 ;
  693 :out2<= 1 ;
  694 :out2<= 1 ;
  695 :out2<= 1 ;
  696 :out2<= 1 ;
  697 :out2<= 1 ;
  698 :out2<= 1 ;
  699 :out2<= 1 ;
  700 :out2<= 1 ;
  701 :out2<= 1 ;
  702 :out2<= 1 ;
  703 :out2<= 1 ;
  704 :out2<= 0 ;
  705 :out2<= 0 ;
  706 :out2<= 0 ;
  707 :out2<= 1 ;
  708 :out2<= 0 ;
  709 :out2<= 1 ;
  710 :out2<= 1 ;
  711 :out2<= 1 ;
  712 :out2<= 0 ;
  713 :out2<= 1 ;
  714 :out2<= 1 ;
  715 :out2<= 1 ;
  716 :out2<= 1 ;
  717 :out2<= 1 ;
  718 :out2<= 1 ;
  719 :out2<= 1 ;
  720 :out2<= 1 ;
  721 :out2<= 1 ;
  722 :out2<= 1 ;
  723 :out2<= 1 ;
  724 :out2<= 1 ;
  725 :out2<= 1 ;
  726 :out2<= 1 ;
  727 :out2<= 1 ;
  728 :out2<= 1 ;
  729 :out2<= 1 ;
  730 :out2<= 1 ;
  731 :out2<= 1 ;
  732 :out2<= 1 ;
  733 :out2<= 1 ;
  734 :out2<= 1 ;
  735 :out2<= 1 ;
  736 :out2<= 1 ;
  737 :out2<= 1 ;
  738 :out2<= 1 ;
  739 :out2<= 1 ;
  740 :out2<= 1 ;
  741 :out2<= 1 ;
  742 :out2<= 1 ;
  743 :out2<= 1 ;
  744 :out2<= 1 ;
  745 :out2<= 1 ;
  746 :out2<= 1 ;
  747 :out2<= 1 ;
  748 :out2<= 1 ;
  749 :out2<= 1 ;
  750 :out2<= 1 ;
  751 :out2<= 1 ;
  752 :out2<= 1 ;
  753 :out2<= 1 ;
  754 :out2<= 1 ;
  755 :out2<= 1 ;
  756 :out2<= 1 ;
  757 :out2<= 1 ;
  758 :out2<= 1 ;
  759 :out2<= 1 ;
  760 :out2<= 1 ;
  761 :out2<= 1 ;
  762 :out2<= 1 ;
  763 :out2<= 1 ;
  764 :out2<= 1 ;
  765 :out2<= 1 ;
  766 :out2<= 1 ;
  767 :out2<= 1 ;
  768 :out2<= 0 ;
  769 :out2<= 0 ;
  770 :out2<= 0 ;
  771 :out2<= 0 ;
  772 :out2<= 0 ;
  773 :out2<= 0 ;
  774 :out2<= 0 ;
  775 :out2<= 1 ;
  776 :out2<= 0 ;
  777 :out2<= 0 ;
  778 :out2<= 0 ;
  779 :out2<= 1 ;
  780 :out2<= 0 ;
  781 :out2<= 1 ;
  782 :out2<= 1 ;
  783 :out2<= 1 ;
  784 :out2<= 0 ;
  785 :out2<= 0 ;
  786 :out2<= 0 ;
  787 :out2<= 1 ;
  788 :out2<= 0 ;
  789 :out2<= 1 ;
  790 :out2<= 1 ;
  791 :out2<= 1 ;
  792 :out2<= 0 ;
  793 :out2<= 1 ;
  794 :out2<= 1 ;
  795 :out2<= 1 ;
  796 :out2<= 1 ;
  797 :out2<= 1 ;
  798 :out2<= 1 ;
  799 :out2<= 1 ;
  800 :out2<= 0 ;
  801 :out2<= 0 ;
  802 :out2<= 0 ;
  803 :out2<= 1 ;
  804 :out2<= 1 ;
  805 :out2<= 1 ;
  806 :out2<= 1 ;
  807 :out2<= 1 ;
  808 :out2<= 1 ;
  809 :out2<= 1 ;
  810 :out2<= 1 ;
  811 :out2<= 1 ;
  812 :out2<= 1 ;
  813 :out2<= 1 ;
  814 :out2<= 1 ;
  815 :out2<= 1 ;
  816 :out2<= 1 ;
  817 :out2<= 1 ;
  818 :out2<= 1 ;
  819 :out2<= 1 ;
  820 :out2<= 1 ;
  821 :out2<= 1 ;
  822 :out2<= 1 ;
  823 :out2<= 1 ;
  824 :out2<= 1 ;
  825 :out2<= 1 ;
  826 :out2<= 1 ;
  827 :out2<= 1 ;
  828 :out2<= 1 ;
  829 :out2<= 1 ;
  830 :out2<= 1 ;
  831 :out2<= 1 ;
  832 :out2<= 0 ;
  833 :out2<= 0 ;
  834 :out2<= 1 ;
  835 :out2<= 1 ;
  836 :out2<= 1 ;
  837 :out2<= 1 ;
  838 :out2<= 1 ;
  839 :out2<= 1 ;
  840 :out2<= 1 ;
  841 :out2<= 1 ;
  842 :out2<= 1 ;
  843 :out2<= 1 ;
  844 :out2<= 1 ;
  845 :out2<= 1 ;
  846 :out2<= 1 ;
  847 :out2<= 1 ;
  848 :out2<= 1 ;
  849 :out2<= 1 ;
  850 :out2<= 1 ;
  851 :out2<= 1 ;
  852 :out2<= 1 ;
  853 :out2<= 1 ;
  854 :out2<= 1 ;
  855 :out2<= 1 ;
  856 :out2<= 1 ;
  857 :out2<= 1 ;
  858 :out2<= 1 ;
  859 :out2<= 1 ;
  860 :out2<= 1 ;
  861 :out2<= 1 ;
  862 :out2<= 1 ;
  863 :out2<= 1 ;
  864 :out2<= 1 ;
  865 :out2<= 1 ;
  866 :out2<= 1 ;
  867 :out2<= 1 ;
  868 :out2<= 1 ;
  869 :out2<= 1 ;
  870 :out2<= 1 ;
  871 :out2<= 1 ;
  872 :out2<= 1 ;
  873 :out2<= 1 ;
  874 :out2<= 1 ;
  875 :out2<= 1 ;
  876 :out2<= 1 ;
  877 :out2<= 1 ;
  878 :out2<= 1 ;
  879 :out2<= 1 ;
  880 :out2<= 1 ;
  881 :out2<= 1 ;
  882 :out2<= 1 ;
  883 :out2<= 1 ;
  884 :out2<= 1 ;
  885 :out2<= 1 ;
  886 :out2<= 1 ;
  887 :out2<= 1 ;
  888 :out2<= 1 ;
  889 :out2<= 1 ;
  890 :out2<= 1 ;
  891 :out2<= 1 ;
  892 :out2<= 1 ;
  893 :out2<= 1 ;
  894 :out2<= 1 ;
  895 :out2<= 1 ;
  896 :out2<= 0 ;
  897 :out2<= 1 ;
  898 :out2<= 1 ;
  899 :out2<= 1 ;
  900 :out2<= 1 ;
  901 :out2<= 1 ;
  902 :out2<= 1 ;
  903 :out2<= 1 ;
  904 :out2<= 1 ;
  905 :out2<= 1 ;
  906 :out2<= 1 ;
  907 :out2<= 1 ;
  908 :out2<= 1 ;
  909 :out2<= 1 ;
  910 :out2<= 1 ;
  911 :out2<= 1 ;
  912 :out2<= 1 ;
  913 :out2<= 1 ;
  914 :out2<= 1 ;
  915 :out2<= 1 ;
  916 :out2<= 1 ;
  917 :out2<= 1 ;
  918 :out2<= 1 ;
  919 :out2<= 1 ;
  920 :out2<= 1 ;
  921 :out2<= 1 ;
  922 :out2<= 1 ;
  923 :out2<= 1 ;
  924 :out2<= 1 ;
  925 :out2<= 1 ;
  926 :out2<= 1 ;
  927 :out2<= 1 ;
  928 :out2<= 1 ;
  929 :out2<= 1 ;
  930 :out2<= 1 ;
  931 :out2<= 1 ;
  932 :out2<= 1 ;
  933 :out2<= 1 ;
  934 :out2<= 1 ;
  935 :out2<= 1 ;
  936 :out2<= 1 ;
  937 :out2<= 1 ;
  938 :out2<= 1 ;
  939 :out2<= 1 ;
  940 :out2<= 1 ;
  941 :out2<= 1 ;
  942 :out2<= 1 ;
  943 :out2<= 1 ;
  944 :out2<= 1 ;
  945 :out2<= 1 ;
  946 :out2<= 1 ;
  947 :out2<= 1 ;
  948 :out2<= 1 ;
  949 :out2<= 1 ;
  950 :out2<= 1 ;
  951 :out2<= 1 ;
  952 :out2<= 1 ;
  953 :out2<= 1 ;
  954 :out2<= 1 ;
  955 :out2<= 1 ;
  956 :out2<= 1 ;
  957 :out2<= 1 ;
  958 :out2<= 1 ;
  959 :out2<= 1 ;
  960 :out2<= 1 ;
  961 :out2<= 1 ;
  962 :out2<= 1 ;
  963 :out2<= 1 ;
  964 :out2<= 1 ;
  965 :out2<= 1 ;
  966 :out2<= 1 ;
  967 :out2<= 1 ;
  968 :out2<= 1 ;
  969 :out2<= 1 ;
  970 :out2<= 1 ;
  971 :out2<= 1 ;
  972 :out2<= 1 ;
  973 :out2<= 1 ;
  974 :out2<= 1 ;
  975 :out2<= 1 ;
  976 :out2<= 1 ;
  977 :out2<= 1 ;
  978 :out2<= 1 ;
  979 :out2<= 1 ;
  980 :out2<= 1 ;
  981 :out2<= 1 ;
  982 :out2<= 1 ;
  983 :out2<= 1 ;
  984 :out2<= 1 ;
  985 :out2<= 1 ;
  986 :out2<= 1 ;
  987 :out2<= 1 ;
  988 :out2<= 1 ;
  989 :out2<= 1 ;
  990 :out2<= 1 ;
  991 :out2<= 1 ;
  992 :out2<= 1 ;
  993 :out2<= 1 ;
  994 :out2<= 1 ;
  995 :out2<= 1 ;
  996 :out2<= 1 ;
  997 :out2<= 1 ;
  998 :out2<= 1 ;
  999 :out2<= 1 ;
  1000 :out2<= 1 ;
  1001 :out2<= 1 ;
  1002 :out2<= 1 ;
  1003 :out2<= 1 ;
  1004 :out2<= 1 ;
  1005 :out2<= 1 ;
  1006 :out2<= 1 ;
  1007 :out2<= 1 ;
  1008 :out2<= 1 ;
  1009 :out2<= 1 ;
  1010 :out2<= 1 ;
  1011 :out2<= 1 ;
  1012 :out2<= 1 ;
  1013 :out2<= 1 ;
  1014 :out2<= 1 ;
  1015 :out2<= 1 ;
  1016 :out2<= 1 ;
  1017 :out2<= 1 ;
  1018 :out2<= 1 ;
  1019 :out2<= 1 ;
  1020 :out2<= 1 ;
  1021 :out2<= 1 ;
  1022 :out2<= 1 ;
  1023 :out2<= 1 ;
 endcase
end

else begin
  out <= 0;
  out2 <= 0;
end

end
endmodule


