module opcode #(parameter P = 128) (clk, rst, channel, I_program_counter,O_opcode, O_opcode_next, O_opcode_delay,
        O_Nv,O_Nv_next, O_part_count,O_part_count_next, O_address, O_address_next, O_opcode_before, O_Nv_before, O_bit_count);
        input clk,rst;
        input channel;
        input [15:0] I_program_counter;
        output [3:0] O_opcode,O_opcode_next, O_opcode_before, O_opcode_delay;
        output [10:0] O_Nv, O_Nv_next, O_Nv_before;
        output [3:0] O_part_count, O_part_count_next;
        output [9:0] O_address, O_address_next;
        output [12:0] O_bit_count;
        localparam TYPE1     = 4'b0000;
        localparam TYPE2     = 4'b0001;
        localparam BOTTOM    = 4'b0010;
        localparam TYPE3     = 4'b0011;
        localparam IDLE      = 4'b1011;

        reg [3:0] L_opcode, L_opcode_next, L_opcode_before, L_opcode_delay;
        reg [10:0] L_Nv,L_Nv_next,L_Nv_before, L_Nv_delay;
        reg [3:0] L_part_count, L_part_count_next, L_part_count_delay;
        reg [9:0] Address, Address_next, Address_delay;
        reg[12:0] L_bit_count;
        
        // assignment of outputs
        assign O_opcode = L_opcode;
        assign O_opcode_delay = L_opcode_delay;
        assign O_opcode_next = L_opcode_next;
        assign O_opcode_before = L_opcode_before;
        assign O_Nv = L_Nv;
        assign O_Nv_next = L_Nv_next;
        assign O_Nv_before = L_Nv_before;
        assign O_part_count = L_part_count;
        assign O_part_count_next = L_part_count_next;
        assign O_address = Address;
        assign O_address_next = Address_next;
        assign O_bit_count = L_bit_count;


        wire islast, oprand;
       assign islast = (L_Nv_next) > (2*P*(1+L_part_count_next));
       assign oprand = (L_opcode_next==TYPE1||L_opcode_next==TYPE2);

       always @(posedge clk)
     begin       
           if(!rst) begin
                L_Nv_before <= L_Nv;        
                L_Nv <= L_Nv_delay;
                L_Nv_delay <= L_Nv_next;

                L_opcode_before <= L_opcode;
                L_opcode <= L_opcode_delay;
                L_opcode_delay <= L_opcode_next;


                L_part_count <= L_part_count_delay;
                L_part_count_delay <= L_part_count_next;

//                Address_before <= Address;       
                L_bit_count <= (L_bit_count+2*(L_opcode==BOTTOM));

                Address <= Address_delay;
                Address_delay <= Address_next;
            end
            else begin
              L_bit_count <= 0;
              L_Nv                          <=1024; 
              L_Nv_before                          <=1024; 
              L_Nv_delay                          <=1024; 

              L_opcode_before <= TYPE1;
              L_opcode <= TYPE1;
              L_opcode_delay <= TYPE1;


              L_part_count <= 0;
              L_part_count_delay <= 0;

              Address <= 0;
              Address_delay <= 0;
            end
        end



        always @(posedge clk) begin
            if(rst) begin
            
            L_Nv_next                     <=1024;
            L_opcode_next <= TYPE1;
            L_part_count_next <= 0;
            // Address <= -1;
            Address_next <= 0;
            end
            else begin
           if (channel) begin
              case (L_Nv_next)
                1024 : L_Nv_next <= islast ? 1024 : 512;
                512 : L_Nv_next <= islast ?  512 : (oprand?256:1024);
                256 : L_Nv_next <= islast ? 256 : (oprand?128:512);
                128 : L_Nv_next <= oprand ? 64 : 256;
                64 : L_Nv_next <= oprand ? 32 : 128;
                32 : L_Nv_next <= oprand ? 16 : 64;
                16 : L_Nv_next <= oprand ? 8 : 32;
                8 : L_Nv_next <= oprand ? 4 : 16;
                4 : L_Nv_next <= oprand ? 2 : 8;
                2 : L_Nv_next <= 4;
                default: L_Nv_next <= 1024;
              endcase

              case (L_opcode_next)
                TYPE1 : L_opcode_next <= islast ? TYPE1 : ( (L_Nv_next==4) ? BOTTOM : TYPE1 );
                TYPE2 : L_opcode_next <= islast ? TYPE2 : ( (L_Nv_next==4) ? BOTTOM : TYPE1 );
                TYPE3 : L_opcode_next <= islast ? TYPE3 : ( (Address_next[0]) ? TYPE3 : TYPE2);
                BOTTOM : L_opcode_next <= Address_next[0] ? TYPE3 : TYPE2 ;
                default: L_opcode_next <= TYPE1;
              endcase

                case (L_part_count_next)
                  0 : L_part_count_next <= (L_Nv_next>2*P) ? 1 : 0;
                  1 : L_part_count_next <= (L_Nv_next>4*P) ? 2 : 0;
                  2 : L_part_count_next <= (L_Nv_next>4*P) ? 3 : 0;
                  3 : L_part_count_next <=  0;
                  // 4 : L_part_count_next <= (L_Nv_next>8*P) ? 5 : 0;
                  // 5 : L_part_count_next <= (L_Nv_next>8*P) ? 6 : 0;
                  // 6 : L_part_count_next <= (L_Nv_next>8*P) ? 7 : 0;
                  // 7 : L_part_count_next <= 0;
                  default: L_part_count_next <= 0;
                endcase


          



       case(I_program_counter)
          9 : Address_next<= 1 ;
          12 : Address_next<= 1 ;
          13 : Address_next<= 2 ;
          15 : Address_next<= 3 ;
          16 : Address_next<= 1 ;
          19 : Address_next<= 1 ;
          20 : Address_next<= 2 ;
          21 : Address_next<= 4 ;
          23 : Address_next<= 5 ;
          24 : Address_next<= 2 ;
          26 : Address_next<= 3 ;
          27 : Address_next<= 6 ;
          29 : Address_next<= 7 ;
          30 : Address_next<= 3 ;
          31 : Address_next<= 1 ;
          34 : Address_next<= 1 ;
          35 : Address_next<= 2 ;
          36 : Address_next<= 4 ;
          37 : Address_next<= 8 ;
          39 : Address_next<= 9 ;
          40 : Address_next<= 4 ;
          42 : Address_next<= 5 ;
          43 : Address_next<= 10 ;
          45 : Address_next<= 11 ;
          46 : Address_next<= 5 ;
          47 : Address_next<= 2 ;
          49 : Address_next<= 3 ;
          50 : Address_next<= 6 ;
          51 : Address_next<= 12 ;
          53 : Address_next<= 13 ;
          54 : Address_next<= 6 ;
          56 : Address_next<= 7 ;
          57 : Address_next<= 14 ;
          59 : Address_next<= 15 ;
          60 : Address_next<= 7 ;
          61 : Address_next<= 3 ;
          62 : Address_next<= 1 ;
          65 : Address_next<= 1 ;
          66 : Address_next<= 2 ;
          67 : Address_next<= 4 ;
          68 : Address_next<= 8 ;
          69 : Address_next<= 16 ;
          71 : Address_next<= 17 ;
          72 : Address_next<= 8 ;
          74 : Address_next<= 9 ;
          75 : Address_next<= 18 ;
          77 : Address_next<= 19 ;
          78 : Address_next<= 9 ;
          79 : Address_next<= 4 ;
          81 : Address_next<= 5 ;
          82 : Address_next<= 10 ;
          83 : Address_next<= 20 ;
          85 : Address_next<= 21 ;
          86 : Address_next<= 10 ;
          88 : Address_next<= 11 ;
          89 : Address_next<= 22 ;
          91 : Address_next<= 23 ;
          92 : Address_next<= 11 ;
          93 : Address_next<= 5 ;
          94 : Address_next<= 2 ;
          96 : Address_next<= 3 ;
          97 : Address_next<= 6 ;
          98 : Address_next<= 12 ;
          99 : Address_next<= 24 ;
          101 : Address_next<= 25 ;
          102 : Address_next<= 12 ;
          104 : Address_next<= 13 ;
          105 : Address_next<= 26 ;
          107 : Address_next<= 27 ;
          108 : Address_next<= 13 ;
          109 : Address_next<= 6 ;
          111 : Address_next<= 7 ;
          112 : Address_next<= 14 ;
          113 : Address_next<= 28 ;
          115 : Address_next<= 29 ;
          116 : Address_next<= 14 ;
          118 : Address_next<= 15 ;
          119 : Address_next<= 30 ;
          121 : Address_next<= 31 ;
          122 : Address_next<= 15 ;
          123 : Address_next<= 7 ;
          124 : Address_next<= 3 ;
          125 : Address_next<= 1 ;
          128 : Address_next<= 1 ;
          129 : Address_next<= 2 ;
          130 : Address_next<= 4 ;
          131 : Address_next<= 8 ;
          132 : Address_next<= 16 ;
          133 : Address_next<= 32 ;
          135 : Address_next<= 33 ;
          136 : Address_next<= 16 ;
          138 : Address_next<= 17 ;
          139 : Address_next<= 34 ;
          141 : Address_next<= 35 ;
          142 : Address_next<= 17 ;
          143 : Address_next<= 8 ;
          145 : Address_next<= 9 ;
          146 : Address_next<= 18 ;
          147 : Address_next<= 36 ;
          149 : Address_next<= 37 ;
          150 : Address_next<= 18 ;
          152 : Address_next<= 19 ;
          153 : Address_next<= 38 ;
          155 : Address_next<= 39 ;
          156 : Address_next<= 19 ;
          157 : Address_next<= 9 ;
          158 : Address_next<= 4 ;
          160 : Address_next<= 5 ;
          161 : Address_next<= 10 ;
          162 : Address_next<= 20 ;
          163 : Address_next<= 40 ;
          165 : Address_next<= 41 ;
          166 : Address_next<= 20 ;
          168 : Address_next<= 21 ;
          169 : Address_next<= 42 ;
          171 : Address_next<= 43 ;
          172 : Address_next<= 21 ;
          173 : Address_next<= 10 ;
          175 : Address_next<= 11 ;
          176 : Address_next<= 22 ;
          177 : Address_next<= 44 ;
          179 : Address_next<= 45 ;
          180 : Address_next<= 22 ;
          182 : Address_next<= 23 ;
          183 : Address_next<= 46 ;
          185 : Address_next<= 47 ;
          186 : Address_next<= 23 ;
          187 : Address_next<= 11 ;
          188 : Address_next<= 5 ;
          189 : Address_next<= 2 ;
          191 : Address_next<= 3 ;
          192 : Address_next<= 6 ;
          193 : Address_next<= 12 ;
          194 : Address_next<= 24 ;
          195 : Address_next<= 48 ;
          197 : Address_next<= 49 ;
          198 : Address_next<= 24 ;
          200 : Address_next<= 25 ;
          201 : Address_next<= 50 ;
          203 : Address_next<= 51 ;
          204 : Address_next<= 25 ;
          205 : Address_next<= 12 ;
          207 : Address_next<= 13 ;
          208 : Address_next<= 26 ;
          209 : Address_next<= 52 ;
          211 : Address_next<= 53 ;
          212 : Address_next<= 26 ;
          214 : Address_next<= 27 ;
          215 : Address_next<= 54 ;
          217 : Address_next<= 55 ;
          218 : Address_next<= 27 ;
          219 : Address_next<= 13 ;
          220 : Address_next<= 6 ;
          222 : Address_next<= 7 ;
          223 : Address_next<= 14 ;
          224 : Address_next<= 28 ;
          225 : Address_next<= 56 ;
          227 : Address_next<= 57 ;
          228 : Address_next<= 28 ;
          230 : Address_next<= 29 ;
          231 : Address_next<= 58 ;
          233 : Address_next<= 59 ;
          234 : Address_next<= 29 ;
          235 : Address_next<= 14 ;
          237 : Address_next<= 15 ;
          238 : Address_next<= 30 ;
          239 : Address_next<= 60 ;
          241 : Address_next<= 61 ;
          242 : Address_next<= 30 ;
          244 : Address_next<= 31 ;
          245 : Address_next<= 62 ;
          247 : Address_next<= 63 ;
          248 : Address_next<= 31 ;
          249 : Address_next<= 15 ;
          250 : Address_next<= 7 ;
          251 : Address_next<= 3 ;
          252 : Address_next<= 1 ;
          255 : Address_next<= 1 ;
          256 : Address_next<= 2 ;
          257 : Address_next<= 4 ;
          258 : Address_next<= 8 ;
          259 : Address_next<= 16 ;
          260 : Address_next<= 32 ;
          261 : Address_next<= 64 ;
          263 : Address_next<= 65 ;
          264 : Address_next<= 32 ;
          266 : Address_next<= 33 ;
          267 : Address_next<= 66 ;
          269 : Address_next<= 67 ;
          270 : Address_next<= 33 ;
          271 : Address_next<= 16 ;
          273 : Address_next<= 17 ;
          274 : Address_next<= 34 ;
          275 : Address_next<= 68 ;
          277 : Address_next<= 69 ;
          278 : Address_next<= 34 ;
          280 : Address_next<= 35 ;
          281 : Address_next<= 70 ;
          283 : Address_next<= 71 ;
          284 : Address_next<= 35 ;
          285 : Address_next<= 17 ;
          286 : Address_next<= 8 ;
          288 : Address_next<= 9 ;
          289 : Address_next<= 18 ;
          290 : Address_next<= 36 ;
          291 : Address_next<= 72 ;
          293 : Address_next<= 73 ;
          294 : Address_next<= 36 ;
          296 : Address_next<= 37 ;
          297 : Address_next<= 74 ;
          299 : Address_next<= 75 ;
          300 : Address_next<= 37 ;
          301 : Address_next<= 18 ;
          303 : Address_next<= 19 ;
          304 : Address_next<= 38 ;
          305 : Address_next<= 76 ;
          307 : Address_next<= 77 ;
          308 : Address_next<= 38 ;
          310 : Address_next<= 39 ;
          311 : Address_next<= 78 ;
          313 : Address_next<= 79 ;
          314 : Address_next<= 39 ;
          315 : Address_next<= 19 ;
          316 : Address_next<= 9 ;
          317 : Address_next<= 4 ;
          319 : Address_next<= 5 ;
          320 : Address_next<= 10 ;
          321 : Address_next<= 20 ;
          322 : Address_next<= 40 ;
          323 : Address_next<= 80 ;
          325 : Address_next<= 81 ;
          326 : Address_next<= 40 ;
          328 : Address_next<= 41 ;
          329 : Address_next<= 82 ;
          331 : Address_next<= 83 ;
          332 : Address_next<= 41 ;
          333 : Address_next<= 20 ;
          335 : Address_next<= 21 ;
          336 : Address_next<= 42 ;
          337 : Address_next<= 84 ;
          339 : Address_next<= 85 ;
          340 : Address_next<= 42 ;
          342 : Address_next<= 43 ;
          343 : Address_next<= 86 ;
          345 : Address_next<= 87 ;
          346 : Address_next<= 43 ;
          347 : Address_next<= 21 ;
          348 : Address_next<= 10 ;
          350 : Address_next<= 11 ;
          351 : Address_next<= 22 ;
          352 : Address_next<= 44 ;
          353 : Address_next<= 88 ;
          355 : Address_next<= 89 ;
          356 : Address_next<= 44 ;
          358 : Address_next<= 45 ;
          359 : Address_next<= 90 ;
          361 : Address_next<= 91 ;
          362 : Address_next<= 45 ;
          363 : Address_next<= 22 ;
          365 : Address_next<= 23 ;
          366 : Address_next<= 46 ;
          367 : Address_next<= 92 ;
          369 : Address_next<= 93 ;
          370 : Address_next<= 46 ;
          372 : Address_next<= 47 ;
          373 : Address_next<= 94 ;
          375 : Address_next<= 95 ;
          376 : Address_next<= 47 ;
          377 : Address_next<= 23 ;
          378 : Address_next<= 11 ;
          379 : Address_next<= 5 ;
          380 : Address_next<= 2 ;
          382 : Address_next<= 3 ;
          383 : Address_next<= 6 ;
          384 : Address_next<= 12 ;
          385 : Address_next<= 24 ;
          386 : Address_next<= 48 ;
          387 : Address_next<= 96 ;
          389 : Address_next<= 97 ;
          390 : Address_next<= 48 ;
          392 : Address_next<= 49 ;
          393 : Address_next<= 98 ;
          395 : Address_next<= 99 ;
          396 : Address_next<= 49 ;
          397 : Address_next<= 24 ;
          399 : Address_next<= 25 ;
          400 : Address_next<= 50 ;
          401 : Address_next<= 100 ;
          403 : Address_next<= 101 ;
          404 : Address_next<= 50 ;
          406 : Address_next<= 51 ;
          407 : Address_next<= 102 ;
          409 : Address_next<= 103 ;
          410 : Address_next<= 51 ;
          411 : Address_next<= 25 ;
          412 : Address_next<= 12 ;
          414 : Address_next<= 13 ;
          415 : Address_next<= 26 ;
          416 : Address_next<= 52 ;
          417 : Address_next<= 104 ;
          419 : Address_next<= 105 ;
          420 : Address_next<= 52 ;
          422 : Address_next<= 53 ;
          423 : Address_next<= 106 ;
          425 : Address_next<= 107 ;
          426 : Address_next<= 53 ;
          427 : Address_next<= 26 ;
          429 : Address_next<= 27 ;
          430 : Address_next<= 54 ;
          431 : Address_next<= 108 ;
          433 : Address_next<= 109 ;
          434 : Address_next<= 54 ;
          436 : Address_next<= 55 ;
          437 : Address_next<= 110 ;
          439 : Address_next<= 111 ;
          440 : Address_next<= 55 ;
          441 : Address_next<= 27 ;
          442 : Address_next<= 13 ;
          443 : Address_next<= 6 ;
          445 : Address_next<= 7 ;
          446 : Address_next<= 14 ;
          447 : Address_next<= 28 ;
          448 : Address_next<= 56 ;
          449 : Address_next<= 112 ;
          451 : Address_next<= 113 ;
          452 : Address_next<= 56 ;
          454 : Address_next<= 57 ;
          455 : Address_next<= 114 ;
          457 : Address_next<= 115 ;
          458 : Address_next<= 57 ;
          459 : Address_next<= 28 ;
          461 : Address_next<= 29 ;
          462 : Address_next<= 58 ;
          463 : Address_next<= 116 ;
          465 : Address_next<= 117 ;
          466 : Address_next<= 58 ;
          468 : Address_next<= 59 ;
          469 : Address_next<= 118 ;
          471 : Address_next<= 119 ;
          472 : Address_next<= 59 ;
          473 : Address_next<= 29 ;
          474 : Address_next<= 14 ;
          476 : Address_next<= 15 ;
          477 : Address_next<= 30 ;
          478 : Address_next<= 60 ;
          479 : Address_next<= 120 ;
          481 : Address_next<= 121 ;
          482 : Address_next<= 60 ;
          484 : Address_next<= 61 ;
          485 : Address_next<= 122 ;
          487 : Address_next<= 123 ;
          488 : Address_next<= 61 ;
          489 : Address_next<= 30 ;
          491 : Address_next<= 31 ;
          492 : Address_next<= 62 ;
          493 : Address_next<= 124 ;
          495 : Address_next<= 125 ;
          496 : Address_next<= 62 ;
          498 : Address_next<= 63 ;
          499 : Address_next<= 126 ;
          501 : Address_next<= 127 ;
          502 : Address_next<= 63 ;
          503 : Address_next<= 31 ;
          504 : Address_next<= 15 ;
          505 : Address_next<= 7 ;
          506 : Address_next<= 3 ;
          507 : Address_next<= 1 ;
          510 : Address_next<= 1 ;
          511 : Address_next<= 2 ;
          512 : Address_next<= 4 ;
          513 : Address_next<= 8 ;
          514 : Address_next<= 16 ;
          515 : Address_next<= 32 ;
          516 : Address_next<= 64 ;
          517 : Address_next<= 128 ;
          519 : Address_next<= 129 ;
          520 : Address_next<= 64 ;
          522 : Address_next<= 65 ;
          523 : Address_next<= 130 ;
          525 : Address_next<= 131 ;
          526 : Address_next<= 65 ;
          527 : Address_next<= 32 ;
          529 : Address_next<= 33 ;
          530 : Address_next<= 66 ;
          531 : Address_next<= 132 ;
          533 : Address_next<= 133 ;
          534 : Address_next<= 66 ;
          536 : Address_next<= 67 ;
          537 : Address_next<= 134 ;
          539 : Address_next<= 135 ;
          540 : Address_next<= 67 ;
          541 : Address_next<= 33 ;
          542 : Address_next<= 16 ;
          544 : Address_next<= 17 ;
          545 : Address_next<= 34 ;
          546 : Address_next<= 68 ;
          547 : Address_next<= 136 ;
          549 : Address_next<= 137 ;
          550 : Address_next<= 68 ;
          552 : Address_next<= 69 ;
          553 : Address_next<= 138 ;
          555 : Address_next<= 139 ;
          556 : Address_next<= 69 ;
          557 : Address_next<= 34 ;
          559 : Address_next<= 35 ;
          560 : Address_next<= 70 ;
          561 : Address_next<= 140 ;
          563 : Address_next<= 141 ;
          564 : Address_next<= 70 ;
          566 : Address_next<= 71 ;
          567 : Address_next<= 142 ;
          569 : Address_next<= 143 ;
          570 : Address_next<= 71 ;
          571 : Address_next<= 35 ;
          572 : Address_next<= 17 ;
          573 : Address_next<= 8 ;
          575 : Address_next<= 9 ;
          576 : Address_next<= 18 ;
          577 : Address_next<= 36 ;
          578 : Address_next<= 72 ;
          579 : Address_next<= 144 ;
          581 : Address_next<= 145 ;
          582 : Address_next<= 72 ;
          584 : Address_next<= 73 ;
          585 : Address_next<= 146 ;
          587 : Address_next<= 147 ;
          588 : Address_next<= 73 ;
          589 : Address_next<= 36 ;
          591 : Address_next<= 37 ;
          592 : Address_next<= 74 ;
          593 : Address_next<= 148 ;
          595 : Address_next<= 149 ;
          596 : Address_next<= 74 ;
          598 : Address_next<= 75 ;
          599 : Address_next<= 150 ;
          601 : Address_next<= 151 ;
          602 : Address_next<= 75 ;
          603 : Address_next<= 37 ;
          604 : Address_next<= 18 ;
          606 : Address_next<= 19 ;
          607 : Address_next<= 38 ;
          608 : Address_next<= 76 ;
          609 : Address_next<= 152 ;
          611 : Address_next<= 153 ;
          612 : Address_next<= 76 ;
          614 : Address_next<= 77 ;
          615 : Address_next<= 154 ;
          617 : Address_next<= 155 ;
          618 : Address_next<= 77 ;
          619 : Address_next<= 38 ;
          621 : Address_next<= 39 ;
          622 : Address_next<= 78 ;
          623 : Address_next<= 156 ;
          625 : Address_next<= 157 ;
          626 : Address_next<= 78 ;
          628 : Address_next<= 79 ;
          629 : Address_next<= 158 ;
          631 : Address_next<= 159 ;
          632 : Address_next<= 79 ;
          633 : Address_next<= 39 ;
          634 : Address_next<= 19 ;
          635 : Address_next<= 9 ;
          636 : Address_next<= 4 ;
          638 : Address_next<= 5 ;
          639 : Address_next<= 10 ;
          640 : Address_next<= 20 ;
          641 : Address_next<= 40 ;
          642 : Address_next<= 80 ;
          643 : Address_next<= 160 ;
          645 : Address_next<= 161 ;
          646 : Address_next<= 80 ;
          648 : Address_next<= 81 ;
          649 : Address_next<= 162 ;
          651 : Address_next<= 163 ;
          652 : Address_next<= 81 ;
          653 : Address_next<= 40 ;
          655 : Address_next<= 41 ;
          656 : Address_next<= 82 ;
          657 : Address_next<= 164 ;
          659 : Address_next<= 165 ;
          660 : Address_next<= 82 ;
          662 : Address_next<= 83 ;
          663 : Address_next<= 166 ;
          665 : Address_next<= 167 ;
          666 : Address_next<= 83 ;
          667 : Address_next<= 41 ;
          668 : Address_next<= 20 ;
          670 : Address_next<= 21 ;
          671 : Address_next<= 42 ;
          672 : Address_next<= 84 ;
          673 : Address_next<= 168 ;
          675 : Address_next<= 169 ;
          676 : Address_next<= 84 ;
          678 : Address_next<= 85 ;
          679 : Address_next<= 170 ;
          681 : Address_next<= 171 ;
          682 : Address_next<= 85 ;
          683 : Address_next<= 42 ;
          685 : Address_next<= 43 ;
          686 : Address_next<= 86 ;
          687 : Address_next<= 172 ;
          689 : Address_next<= 173 ;
          690 : Address_next<= 86 ;
          692 : Address_next<= 87 ;
          693 : Address_next<= 174 ;
          695 : Address_next<= 175 ;
          696 : Address_next<= 87 ;
          697 : Address_next<= 43 ;
          698 : Address_next<= 21 ;
          699 : Address_next<= 10 ;
          701 : Address_next<= 11 ;
          702 : Address_next<= 22 ;
          703 : Address_next<= 44 ;
          704 : Address_next<= 88 ;
          705 : Address_next<= 176 ;
          707 : Address_next<= 177 ;
          708 : Address_next<= 88 ;
          710 : Address_next<= 89 ;
          711 : Address_next<= 178 ;
          713 : Address_next<= 179 ;
          714 : Address_next<= 89 ;
          715 : Address_next<= 44 ;
          717 : Address_next<= 45 ;
          718 : Address_next<= 90 ;
          719 : Address_next<= 180 ;
          721 : Address_next<= 181 ;
          722 : Address_next<= 90 ;
          724 : Address_next<= 91 ;
          725 : Address_next<= 182 ;
          727 : Address_next<= 183 ;
          728 : Address_next<= 91 ;
          729 : Address_next<= 45 ;
          730 : Address_next<= 22 ;
          732 : Address_next<= 23 ;
          733 : Address_next<= 46 ;
          734 : Address_next<= 92 ;
          735 : Address_next<= 184 ;
          737 : Address_next<= 185 ;
          738 : Address_next<= 92 ;
          740 : Address_next<= 93 ;
          741 : Address_next<= 186 ;
          743 : Address_next<= 187 ;
          744 : Address_next<= 93 ;
          745 : Address_next<= 46 ;
          747 : Address_next<= 47 ;
          748 : Address_next<= 94 ;
          749 : Address_next<= 188 ;
          751 : Address_next<= 189 ;
          752 : Address_next<= 94 ;
          754 : Address_next<= 95 ;
          755 : Address_next<= 190 ;
          757 : Address_next<= 191 ;
          758 : Address_next<= 95 ;
          759 : Address_next<= 47 ;
          760 : Address_next<= 23 ;
          761 : Address_next<= 11 ;
          762 : Address_next<= 5 ;
          763 : Address_next<= 2 ;
          765 : Address_next<= 3 ;
          766 : Address_next<= 6 ;
          767 : Address_next<= 12 ;
          768 : Address_next<= 24 ;
          769 : Address_next<= 48 ;
          770 : Address_next<= 96 ;
          771 : Address_next<= 192 ;
          773 : Address_next<= 193 ;
          774 : Address_next<= 96 ;
          776 : Address_next<= 97 ;
          777 : Address_next<= 194 ;
          779 : Address_next<= 195 ;
          780 : Address_next<= 97 ;
          781 : Address_next<= 48 ;
          783 : Address_next<= 49 ;
          784 : Address_next<= 98 ;
          785 : Address_next<= 196 ;
          787 : Address_next<= 197 ;
          788 : Address_next<= 98 ;
          790 : Address_next<= 99 ;
          791 : Address_next<= 198 ;
          793 : Address_next<= 199 ;
          794 : Address_next<= 99 ;
          795 : Address_next<= 49 ;
          796 : Address_next<= 24 ;
          798 : Address_next<= 25 ;
          799 : Address_next<= 50 ;
          800 : Address_next<= 100 ;
          801 : Address_next<= 200 ;
          803 : Address_next<= 201 ;
          804 : Address_next<= 100 ;
          806 : Address_next<= 101 ;
          807 : Address_next<= 202 ;
          809 : Address_next<= 203 ;
          810 : Address_next<= 101 ;
          811 : Address_next<= 50 ;
          813 : Address_next<= 51 ;
          814 : Address_next<= 102 ;
          815 : Address_next<= 204 ;
          817 : Address_next<= 205 ;
          818 : Address_next<= 102 ;
          820 : Address_next<= 103 ;
          821 : Address_next<= 206 ;
          823 : Address_next<= 207 ;
          824 : Address_next<= 103 ;
          825 : Address_next<= 51 ;
          826 : Address_next<= 25 ;
          827 : Address_next<= 12 ;
          829 : Address_next<= 13 ;
          830 : Address_next<= 26 ;
          831 : Address_next<= 52 ;
          832 : Address_next<= 104 ;
          833 : Address_next<= 208 ;
          835 : Address_next<= 209 ;
          836 : Address_next<= 104 ;
          838 : Address_next<= 105 ;
          839 : Address_next<= 210 ;
          841 : Address_next<= 211 ;
          842 : Address_next<= 105 ;
          843 : Address_next<= 52 ;
          845 : Address_next<= 53 ;
          846 : Address_next<= 106 ;
          847 : Address_next<= 212 ;
          849 : Address_next<= 213 ;
          850 : Address_next<= 106 ;
          852 : Address_next<= 107 ;
          853 : Address_next<= 214 ;
          855 : Address_next<= 215 ;
          856 : Address_next<= 107 ;
          857 : Address_next<= 53 ;
          858 : Address_next<= 26 ;
          860 : Address_next<= 27 ;
          861 : Address_next<= 54 ;
          862 : Address_next<= 108 ;
          863 : Address_next<= 216 ;
          865 : Address_next<= 217 ;
          866 : Address_next<= 108 ;
          868 : Address_next<= 109 ;
          869 : Address_next<= 218 ;
          871 : Address_next<= 219 ;
          872 : Address_next<= 109 ;
          873 : Address_next<= 54 ;
          875 : Address_next<= 55 ;
          876 : Address_next<= 110 ;
          877 : Address_next<= 220 ;
          879 : Address_next<= 221 ;
          880 : Address_next<= 110 ;
          882 : Address_next<= 111 ;
          883 : Address_next<= 222 ;
          885 : Address_next<= 223 ;
          886 : Address_next<= 111 ;
          887 : Address_next<= 55 ;
          888 : Address_next<= 27 ;
          889 : Address_next<= 13 ;
          890 : Address_next<= 6 ;
          892 : Address_next<= 7 ;
          893 : Address_next<= 14 ;
          894 : Address_next<= 28 ;
          895 : Address_next<= 56 ;
          896 : Address_next<= 112 ;
          897 : Address_next<= 224 ;
          899 : Address_next<= 225 ;
          900 : Address_next<= 112 ;
          902 : Address_next<= 113 ;
          903 : Address_next<= 226 ;
          905 : Address_next<= 227 ;
          906 : Address_next<= 113 ;
          907 : Address_next<= 56 ;
          909 : Address_next<= 57 ;
          910 : Address_next<= 114 ;
          911 : Address_next<= 228 ;
          913 : Address_next<= 229 ;
          914 : Address_next<= 114 ;
          916 : Address_next<= 115 ;
          917 : Address_next<= 230 ;
          919 : Address_next<= 231 ;
          920 : Address_next<= 115 ;
          921 : Address_next<= 57 ;
          922 : Address_next<= 28 ;
          924 : Address_next<= 29 ;
          925 : Address_next<= 58 ;
          926 : Address_next<= 116 ;
          927 : Address_next<= 232 ;
          929 : Address_next<= 233 ;
          930 : Address_next<= 116 ;
          932 : Address_next<= 117 ;
          933 : Address_next<= 234 ;
          935 : Address_next<= 235 ;
          936 : Address_next<= 117 ;
          937 : Address_next<= 58 ;
          939 : Address_next<= 59 ;
          940 : Address_next<= 118 ;
          941 : Address_next<= 236 ;
          943 : Address_next<= 237 ;
          944 : Address_next<= 118 ;
          946 : Address_next<= 119 ;
          947 : Address_next<= 238 ;
          949 : Address_next<= 239 ;
          950 : Address_next<= 119 ;
          951 : Address_next<= 59 ;
          952 : Address_next<= 29 ;
          953 : Address_next<= 14 ;
          955 : Address_next<= 15 ;
          956 : Address_next<= 30 ;
          957 : Address_next<= 60 ;
          958 : Address_next<= 120 ;
          959 : Address_next<= 240 ;
          961 : Address_next<= 241 ;
          962 : Address_next<= 120 ;
          964 : Address_next<= 121 ;
          965 : Address_next<= 242 ;
          967 : Address_next<= 243 ;
          968 : Address_next<= 121 ;
          969 : Address_next<= 60 ;
          971 : Address_next<= 61 ;
          972 : Address_next<= 122 ;
          973 : Address_next<= 244 ;
          975 : Address_next<= 245 ;
          976 : Address_next<= 122 ;
          978 : Address_next<= 123 ;
          979 : Address_next<= 246 ;
          981 : Address_next<= 247 ;
          982 : Address_next<= 123 ;
          983 : Address_next<= 61 ;
          984 : Address_next<= 30 ;
          986 : Address_next<= 31 ;
          987 : Address_next<= 62 ;
          988 : Address_next<= 124 ;
          989 : Address_next<= 248 ;
          991 : Address_next<= 249 ;
          992 : Address_next<= 124 ;
          994 : Address_next<= 125 ;
          995 : Address_next<= 250 ;
          997 : Address_next<= 251 ;
          998 : Address_next<= 125 ;
          999 : Address_next<= 62 ;
          1001 : Address_next<= 63 ;
          1002 : Address_next<= 126 ;
          1003 : Address_next<= 252 ;
          1005 : Address_next<= 253 ;
          1006 : Address_next<= 126 ;
          1008 : Address_next<= 127 ;
          1009 : Address_next<= 254 ;
          1011 : Address_next<= 255 ;
          1012 : Address_next<= 127 ;
          1013 : Address_next<= 63 ;
          1014 : Address_next<= 31 ;
          1015 : Address_next<= 15 ;
          1016 : Address_next<= 7 ;
          1017 : Address_next<= 3 ;
          1018 : Address_next<= 1 ;
          1022 : Address_next<= 1 ;
          1023 : Address_next<= 2 ;
          1024 : Address_next<= 4 ;
          1025 : Address_next<= 8 ;
          1026 : Address_next<= 16 ;
          1027 : Address_next<= 32 ;
          1028 : Address_next<= 64 ;
          1029 : Address_next<= 128 ;
          1030 : Address_next<= 256 ;
          1032 : Address_next<= 257 ;
          1033 : Address_next<= 128 ;
          1035 : Address_next<= 129 ;
          1036 : Address_next<= 258 ;
          1038 : Address_next<= 259 ;
          1039 : Address_next<= 129 ;
          1040 : Address_next<= 64 ;
          1042 : Address_next<= 65 ;
          1043 : Address_next<= 130 ;
          1044 : Address_next<= 260 ;
          1046 : Address_next<= 261 ;
          1047 : Address_next<= 130 ;
          1049 : Address_next<= 131 ;
          1050 : Address_next<= 262 ;
          1052 : Address_next<= 263 ;
          1053 : Address_next<= 131 ;
          1054 : Address_next<= 65 ;
          1055 : Address_next<= 32 ;
          1057 : Address_next<= 33 ;
          1058 : Address_next<= 66 ;
          1059 : Address_next<= 132 ;
          1060 : Address_next<= 264 ;
          1062 : Address_next<= 265 ;
          1063 : Address_next<= 132 ;
          1065 : Address_next<= 133 ;
          1066 : Address_next<= 266 ;
          1068 : Address_next<= 267 ;
          1069 : Address_next<= 133 ;
          1070 : Address_next<= 66 ;
          1072 : Address_next<= 67 ;
          1073 : Address_next<= 134 ;
          1074 : Address_next<= 268 ;
          1076 : Address_next<= 269 ;
          1077 : Address_next<= 134 ;
          1079 : Address_next<= 135 ;
          1080 : Address_next<= 270 ;
          1082 : Address_next<= 271 ;
          1083 : Address_next<= 135 ;
          1084 : Address_next<= 67 ;
          1085 : Address_next<= 33 ;
          1086 : Address_next<= 16 ;
          1088 : Address_next<= 17 ;
          1089 : Address_next<= 34 ;
          1090 : Address_next<= 68 ;
          1091 : Address_next<= 136 ;
          1092 : Address_next<= 272 ;
          1094 : Address_next<= 273 ;
          1095 : Address_next<= 136 ;
          1097 : Address_next<= 137 ;
          1098 : Address_next<= 274 ;
          1100 : Address_next<= 275 ;
          1101 : Address_next<= 137 ;
          1102 : Address_next<= 68 ;
          1104 : Address_next<= 69 ;
          1105 : Address_next<= 138 ;
          1106 : Address_next<= 276 ;
          1108 : Address_next<= 277 ;
          1109 : Address_next<= 138 ;
          1111 : Address_next<= 139 ;
          1112 : Address_next<= 278 ;
          1114 : Address_next<= 279 ;
          1115 : Address_next<= 139 ;
          1116 : Address_next<= 69 ;
          1117 : Address_next<= 34 ;
          1119 : Address_next<= 35 ;
          1120 : Address_next<= 70 ;
          1121 : Address_next<= 140 ;
          1122 : Address_next<= 280 ;
          1124 : Address_next<= 281 ;
          1125 : Address_next<= 140 ;
          1127 : Address_next<= 141 ;
          1128 : Address_next<= 282 ;
          1130 : Address_next<= 283 ;
          1131 : Address_next<= 141 ;
          1132 : Address_next<= 70 ;
          1134 : Address_next<= 71 ;
          1135 : Address_next<= 142 ;
          1136 : Address_next<= 284 ;
          1138 : Address_next<= 285 ;
          1139 : Address_next<= 142 ;
          1141 : Address_next<= 143 ;
          1142 : Address_next<= 286 ;
          1144 : Address_next<= 287 ;
          1145 : Address_next<= 143 ;
          1146 : Address_next<= 71 ;
          1147 : Address_next<= 35 ;
          1148 : Address_next<= 17 ;
          1149 : Address_next<= 8 ;
          1151 : Address_next<= 9 ;
          1152 : Address_next<= 18 ;
          1153 : Address_next<= 36 ;
          1154 : Address_next<= 72 ;
          1155 : Address_next<= 144 ;
          1156 : Address_next<= 288 ;
          1158 : Address_next<= 289 ;
          1159 : Address_next<= 144 ;
          1161 : Address_next<= 145 ;
          1162 : Address_next<= 290 ;
          1164 : Address_next<= 291 ;
          1165 : Address_next<= 145 ;
          1166 : Address_next<= 72 ;
          1168 : Address_next<= 73 ;
          1169 : Address_next<= 146 ;
          1170 : Address_next<= 292 ;
          1172 : Address_next<= 293 ;
          1173 : Address_next<= 146 ;
          1175 : Address_next<= 147 ;
          1176 : Address_next<= 294 ;
          1178 : Address_next<= 295 ;
          1179 : Address_next<= 147 ;
          1180 : Address_next<= 73 ;
          1181 : Address_next<= 36 ;
          1183 : Address_next<= 37 ;
          1184 : Address_next<= 74 ;
          1185 : Address_next<= 148 ;
          1186 : Address_next<= 296 ;
          1188 : Address_next<= 297 ;
          1189 : Address_next<= 148 ;
          1191 : Address_next<= 149 ;
          1192 : Address_next<= 298 ;
          1194 : Address_next<= 299 ;
          1195 : Address_next<= 149 ;
          1196 : Address_next<= 74 ;
          1198 : Address_next<= 75 ;
          1199 : Address_next<= 150 ;
          1200 : Address_next<= 300 ;
          1202 : Address_next<= 301 ;
          1203 : Address_next<= 150 ;
          1205 : Address_next<= 151 ;
          1206 : Address_next<= 302 ;
          1208 : Address_next<= 303 ;
          1209 : Address_next<= 151 ;
          1210 : Address_next<= 75 ;
          1211 : Address_next<= 37 ;
          1212 : Address_next<= 18 ;
          1214 : Address_next<= 19 ;
          1215 : Address_next<= 38 ;
          1216 : Address_next<= 76 ;
          1217 : Address_next<= 152 ;
          1218 : Address_next<= 304 ;
          1220 : Address_next<= 305 ;
          1221 : Address_next<= 152 ;
          1223 : Address_next<= 153 ;
          1224 : Address_next<= 306 ;
          1226 : Address_next<= 307 ;
          1227 : Address_next<= 153 ;
          1228 : Address_next<= 76 ;
          1230 : Address_next<= 77 ;
          1231 : Address_next<= 154 ;
          1232 : Address_next<= 308 ;
          1234 : Address_next<= 309 ;
          1235 : Address_next<= 154 ;
          1237 : Address_next<= 155 ;
          1238 : Address_next<= 310 ;
          1240 : Address_next<= 311 ;
          1241 : Address_next<= 155 ;
          1242 : Address_next<= 77 ;
          1243 : Address_next<= 38 ;
          1245 : Address_next<= 39 ;
          1246 : Address_next<= 78 ;
          1247 : Address_next<= 156 ;
          1248 : Address_next<= 312 ;
          1250 : Address_next<= 313 ;
          1251 : Address_next<= 156 ;
          1253 : Address_next<= 157 ;
          1254 : Address_next<= 314 ;
          1256 : Address_next<= 315 ;
          1257 : Address_next<= 157 ;
          1258 : Address_next<= 78 ;
          1260 : Address_next<= 79 ;
          1261 : Address_next<= 158 ;
          1262 : Address_next<= 316 ;
          1264 : Address_next<= 317 ;
          1265 : Address_next<= 158 ;
          1267 : Address_next<= 159 ;
          1268 : Address_next<= 318 ;
          1270 : Address_next<= 319 ;
          1271 : Address_next<= 159 ;
          1272 : Address_next<= 79 ;
          1273 : Address_next<= 39 ;
          1274 : Address_next<= 19 ;
          1275 : Address_next<= 9 ;
          1276 : Address_next<= 4 ;
          1278 : Address_next<= 5 ;
          1279 : Address_next<= 10 ;
          1280 : Address_next<= 20 ;
          1281 : Address_next<= 40 ;
          1282 : Address_next<= 80 ;
          1283 : Address_next<= 160 ;
          1284 : Address_next<= 320 ;
          1286 : Address_next<= 321 ;
          1287 : Address_next<= 160 ;
          1289 : Address_next<= 161 ;
          1290 : Address_next<= 322 ;
          1292 : Address_next<= 323 ;
          1293 : Address_next<= 161 ;
          1294 : Address_next<= 80 ;
          1296 : Address_next<= 81 ;
          1297 : Address_next<= 162 ;
          1298 : Address_next<= 324 ;
          1300 : Address_next<= 325 ;
          1301 : Address_next<= 162 ;
          1303 : Address_next<= 163 ;
          1304 : Address_next<= 326 ;
          1306 : Address_next<= 327 ;
          1307 : Address_next<= 163 ;
          1308 : Address_next<= 81 ;
          1309 : Address_next<= 40 ;
          1311 : Address_next<= 41 ;
          1312 : Address_next<= 82 ;
          1313 : Address_next<= 164 ;
          1314 : Address_next<= 328 ;
          1316 : Address_next<= 329 ;
          1317 : Address_next<= 164 ;
          1319 : Address_next<= 165 ;
          1320 : Address_next<= 330 ;
          1322 : Address_next<= 331 ;
          1323 : Address_next<= 165 ;
          1324 : Address_next<= 82 ;
          1326 : Address_next<= 83 ;
          1327 : Address_next<= 166 ;
          1328 : Address_next<= 332 ;
          1330 : Address_next<= 333 ;
          1331 : Address_next<= 166 ;
          1333 : Address_next<= 167 ;
          1334 : Address_next<= 334 ;
          1336 : Address_next<= 335 ;
          1337 : Address_next<= 167 ;
          1338 : Address_next<= 83 ;
          1339 : Address_next<= 41 ;
          1340 : Address_next<= 20 ;
          1342 : Address_next<= 21 ;
          1343 : Address_next<= 42 ;
          1344 : Address_next<= 84 ;
          1345 : Address_next<= 168 ;
          1346 : Address_next<= 336 ;
          1348 : Address_next<= 337 ;
          1349 : Address_next<= 168 ;
          1351 : Address_next<= 169 ;
          1352 : Address_next<= 338 ;
          1354 : Address_next<= 339 ;
          1355 : Address_next<= 169 ;
          1356 : Address_next<= 84 ;
          1358 : Address_next<= 85 ;
          1359 : Address_next<= 170 ;
          1360 : Address_next<= 340 ;
          1362 : Address_next<= 341 ;
          1363 : Address_next<= 170 ;
          1365 : Address_next<= 171 ;
          1366 : Address_next<= 342 ;
          1368 : Address_next<= 343 ;
          1369 : Address_next<= 171 ;
          1370 : Address_next<= 85 ;
          1371 : Address_next<= 42 ;
          1373 : Address_next<= 43 ;
          1374 : Address_next<= 86 ;
          1375 : Address_next<= 172 ;
          1376 : Address_next<= 344 ;
          1378 : Address_next<= 345 ;
          1379 : Address_next<= 172 ;
          1381 : Address_next<= 173 ;
          1382 : Address_next<= 346 ;
          1384 : Address_next<= 347 ;
          1385 : Address_next<= 173 ;
          1386 : Address_next<= 86 ;
          1388 : Address_next<= 87 ;
          1389 : Address_next<= 174 ;
          1390 : Address_next<= 348 ;
          1392 : Address_next<= 349 ;
          1393 : Address_next<= 174 ;
          1395 : Address_next<= 175 ;
          1396 : Address_next<= 350 ;
          1398 : Address_next<= 351 ;
          1399 : Address_next<= 175 ;
          1400 : Address_next<= 87 ;
          1401 : Address_next<= 43 ;
          1402 : Address_next<= 21 ;
          1403 : Address_next<= 10 ;
          1405 : Address_next<= 11 ;
          1406 : Address_next<= 22 ;
          1407 : Address_next<= 44 ;
          1408 : Address_next<= 88 ;
          1409 : Address_next<= 176 ;
          1410 : Address_next<= 352 ;
          1412 : Address_next<= 353 ;
          1413 : Address_next<= 176 ;
          1415 : Address_next<= 177 ;
          1416 : Address_next<= 354 ;
          1418 : Address_next<= 355 ;
          1419 : Address_next<= 177 ;
          1420 : Address_next<= 88 ;
          1422 : Address_next<= 89 ;
          1423 : Address_next<= 178 ;
          1424 : Address_next<= 356 ;
          1426 : Address_next<= 357 ;
          1427 : Address_next<= 178 ;
          1429 : Address_next<= 179 ;
          1430 : Address_next<= 358 ;
          1432 : Address_next<= 359 ;
          1433 : Address_next<= 179 ;
          1434 : Address_next<= 89 ;
          1435 : Address_next<= 44 ;
          1437 : Address_next<= 45 ;
          1438 : Address_next<= 90 ;
          1439 : Address_next<= 180 ;
          1440 : Address_next<= 360 ;
          1442 : Address_next<= 361 ;
          1443 : Address_next<= 180 ;
          1445 : Address_next<= 181 ;
          1446 : Address_next<= 362 ;
          1448 : Address_next<= 363 ;
          1449 : Address_next<= 181 ;
          1450 : Address_next<= 90 ;
          1452 : Address_next<= 91 ;
          1453 : Address_next<= 182 ;
          1454 : Address_next<= 364 ;
          1456 : Address_next<= 365 ;
          1457 : Address_next<= 182 ;
          1459 : Address_next<= 183 ;
          1460 : Address_next<= 366 ;
          1462 : Address_next<= 367 ;
          1463 : Address_next<= 183 ;
          1464 : Address_next<= 91 ;
          1465 : Address_next<= 45 ;
          1466 : Address_next<= 22 ;
          1468 : Address_next<= 23 ;
          1469 : Address_next<= 46 ;
          1470 : Address_next<= 92 ;
          1471 : Address_next<= 184 ;
          1472 : Address_next<= 368 ;
          1474 : Address_next<= 369 ;
          1475 : Address_next<= 184 ;
          1477 : Address_next<= 185 ;
          1478 : Address_next<= 370 ;
          1480 : Address_next<= 371 ;
          1481 : Address_next<= 185 ;
          1482 : Address_next<= 92 ;
          1484 : Address_next<= 93 ;
          1485 : Address_next<= 186 ;
          1486 : Address_next<= 372 ;
          1488 : Address_next<= 373 ;
          1489 : Address_next<= 186 ;
          1491 : Address_next<= 187 ;
          1492 : Address_next<= 374 ;
          1494 : Address_next<= 375 ;
          1495 : Address_next<= 187 ;
          1496 : Address_next<= 93 ;
          1497 : Address_next<= 46 ;
          1499 : Address_next<= 47 ;
          1500 : Address_next<= 94 ;
          1501 : Address_next<= 188 ;
          1502 : Address_next<= 376 ;
          1504 : Address_next<= 377 ;
          1505 : Address_next<= 188 ;
          1507 : Address_next<= 189 ;
          1508 : Address_next<= 378 ;
          1510 : Address_next<= 379 ;
          1511 : Address_next<= 189 ;
          1512 : Address_next<= 94 ;
          1514 : Address_next<= 95 ;
          1515 : Address_next<= 190 ;
          1516 : Address_next<= 380 ;
          1518 : Address_next<= 381 ;
          1519 : Address_next<= 190 ;
          1521 : Address_next<= 191 ;
          1522 : Address_next<= 382 ;
          1524 : Address_next<= 383 ;
          1525 : Address_next<= 191 ;
          1526 : Address_next<= 95 ;
          1527 : Address_next<= 47 ;
          1528 : Address_next<= 23 ;
          1529 : Address_next<= 11 ;
          1530 : Address_next<= 5 ;
          1531 : Address_next<= 2 ;
          1533 : Address_next<= 3 ;
          1534 : Address_next<= 6 ;
          1535 : Address_next<= 12 ;
          1536 : Address_next<= 24 ;
          1537 : Address_next<= 48 ;
          1538 : Address_next<= 96 ;
          1539 : Address_next<= 192 ;
          1540 : Address_next<= 384 ;
          1542 : Address_next<= 385 ;
          1543 : Address_next<= 192 ;
          1545 : Address_next<= 193 ;
          1546 : Address_next<= 386 ;
          1548 : Address_next<= 387 ;
          1549 : Address_next<= 193 ;
          1550 : Address_next<= 96 ;
          1552 : Address_next<= 97 ;
          1553 : Address_next<= 194 ;
          1554 : Address_next<= 388 ;
          1556 : Address_next<= 389 ;
          1557 : Address_next<= 194 ;
          1559 : Address_next<= 195 ;
          1560 : Address_next<= 390 ;
          1562 : Address_next<= 391 ;
          1563 : Address_next<= 195 ;
          1564 : Address_next<= 97 ;
          1565 : Address_next<= 48 ;
          1567 : Address_next<= 49 ;
          1568 : Address_next<= 98 ;
          1569 : Address_next<= 196 ;
          1570 : Address_next<= 392 ;
          1572 : Address_next<= 393 ;
          1573 : Address_next<= 196 ;
          1575 : Address_next<= 197 ;
          1576 : Address_next<= 394 ;
          1578 : Address_next<= 395 ;
          1579 : Address_next<= 197 ;
          1580 : Address_next<= 98 ;
          1582 : Address_next<= 99 ;
          1583 : Address_next<= 198 ;
          1584 : Address_next<= 396 ;
          1586 : Address_next<= 397 ;
          1587 : Address_next<= 198 ;
          1589 : Address_next<= 199 ;
          1590 : Address_next<= 398 ;
          1592 : Address_next<= 399 ;
          1593 : Address_next<= 199 ;
          1594 : Address_next<= 99 ;
          1595 : Address_next<= 49 ;
          1596 : Address_next<= 24 ;
          1598 : Address_next<= 25 ;
          1599 : Address_next<= 50 ;
          1600 : Address_next<= 100 ;
          1601 : Address_next<= 200 ;
          1602 : Address_next<= 400 ;
          1604 : Address_next<= 401 ;
          1605 : Address_next<= 200 ;
          1607 : Address_next<= 201 ;
          1608 : Address_next<= 402 ;
          1610 : Address_next<= 403 ;
          1611 : Address_next<= 201 ;
          1612 : Address_next<= 100 ;
          1614 : Address_next<= 101 ;
          1615 : Address_next<= 202 ;
          1616 : Address_next<= 404 ;
          1618 : Address_next<= 405 ;
          1619 : Address_next<= 202 ;
          1621 : Address_next<= 203 ;
          1622 : Address_next<= 406 ;
          1624 : Address_next<= 407 ;
          1625 : Address_next<= 203 ;
          1626 : Address_next<= 101 ;
          1627 : Address_next<= 50 ;
          1629 : Address_next<= 51 ;
          1630 : Address_next<= 102 ;
          1631 : Address_next<= 204 ;
          1632 : Address_next<= 408 ;
          1634 : Address_next<= 409 ;
          1635 : Address_next<= 204 ;
          1637 : Address_next<= 205 ;
          1638 : Address_next<= 410 ;
          1640 : Address_next<= 411 ;
          1641 : Address_next<= 205 ;
          1642 : Address_next<= 102 ;
          1644 : Address_next<= 103 ;
          1645 : Address_next<= 206 ;
          1646 : Address_next<= 412 ;
          1648 : Address_next<= 413 ;
          1649 : Address_next<= 206 ;
          1651 : Address_next<= 207 ;
          1652 : Address_next<= 414 ;
          1654 : Address_next<= 415 ;
          1655 : Address_next<= 207 ;
          1656 : Address_next<= 103 ;
          1657 : Address_next<= 51 ;
          1658 : Address_next<= 25 ;
          1659 : Address_next<= 12 ;
          1661 : Address_next<= 13 ;
          1662 : Address_next<= 26 ;
          1663 : Address_next<= 52 ;
          1664 : Address_next<= 104 ;
          1665 : Address_next<= 208 ;
          1666 : Address_next<= 416 ;
          1668 : Address_next<= 417 ;
          1669 : Address_next<= 208 ;
          1671 : Address_next<= 209 ;
          1672 : Address_next<= 418 ;
          1674 : Address_next<= 419 ;
          1675 : Address_next<= 209 ;
          1676 : Address_next<= 104 ;
          1678 : Address_next<= 105 ;
          1679 : Address_next<= 210 ;
          1680 : Address_next<= 420 ;
          1682 : Address_next<= 421 ;
          1683 : Address_next<= 210 ;
          1685 : Address_next<= 211 ;
          1686 : Address_next<= 422 ;
          1688 : Address_next<= 423 ;
          1689 : Address_next<= 211 ;
          1690 : Address_next<= 105 ;
          1691 : Address_next<= 52 ;
          1693 : Address_next<= 53 ;
          1694 : Address_next<= 106 ;
          1695 : Address_next<= 212 ;
          1696 : Address_next<= 424 ;
          1698 : Address_next<= 425 ;
          1699 : Address_next<= 212 ;
          1701 : Address_next<= 213 ;
          1702 : Address_next<= 426 ;
          1704 : Address_next<= 427 ;
          1705 : Address_next<= 213 ;
          1706 : Address_next<= 106 ;
          1708 : Address_next<= 107 ;
          1709 : Address_next<= 214 ;
          1710 : Address_next<= 428 ;
          1712 : Address_next<= 429 ;
          1713 : Address_next<= 214 ;
          1715 : Address_next<= 215 ;
          1716 : Address_next<= 430 ;
          1718 : Address_next<= 431 ;
          1719 : Address_next<= 215 ;
          1720 : Address_next<= 107 ;
          1721 : Address_next<= 53 ;
          1722 : Address_next<= 26 ;
          1724 : Address_next<= 27 ;
          1725 : Address_next<= 54 ;
          1726 : Address_next<= 108 ;
          1727 : Address_next<= 216 ;
          1728 : Address_next<= 432 ;
          1730 : Address_next<= 433 ;
          1731 : Address_next<= 216 ;
          1733 : Address_next<= 217 ;
          1734 : Address_next<= 434 ;
          1736 : Address_next<= 435 ;
          1737 : Address_next<= 217 ;
          1738 : Address_next<= 108 ;
          1740 : Address_next<= 109 ;
          1741 : Address_next<= 218 ;
          1742 : Address_next<= 436 ;
          1744 : Address_next<= 437 ;
          1745 : Address_next<= 218 ;
          1747 : Address_next<= 219 ;
          1748 : Address_next<= 438 ;
          1750 : Address_next<= 439 ;
          1751 : Address_next<= 219 ;
          1752 : Address_next<= 109 ;
          1753 : Address_next<= 54 ;
          1755 : Address_next<= 55 ;
          1756 : Address_next<= 110 ;
          1757 : Address_next<= 220 ;
          1758 : Address_next<= 440 ;
          1760 : Address_next<= 441 ;
          1761 : Address_next<= 220 ;
          1763 : Address_next<= 221 ;
          1764 : Address_next<= 442 ;
          1766 : Address_next<= 443 ;
          1767 : Address_next<= 221 ;
          1768 : Address_next<= 110 ;
          1770 : Address_next<= 111 ;
          1771 : Address_next<= 222 ;
          1772 : Address_next<= 444 ;
          1774 : Address_next<= 445 ;
          1775 : Address_next<= 222 ;
          1777 : Address_next<= 223 ;
          1778 : Address_next<= 446 ;
          1780 : Address_next<= 447 ;
          1781 : Address_next<= 223 ;
          1782 : Address_next<= 111 ;
          1783 : Address_next<= 55 ;
          1784 : Address_next<= 27 ;
          1785 : Address_next<= 13 ;
          1786 : Address_next<= 6 ;
          1788 : Address_next<= 7 ;
          1789 : Address_next<= 14 ;
          1790 : Address_next<= 28 ;
          1791 : Address_next<= 56 ;
          1792 : Address_next<= 112 ;
          1793 : Address_next<= 224 ;
          1794 : Address_next<= 448 ;
          1796 : Address_next<= 449 ;
          1797 : Address_next<= 224 ;
          1799 : Address_next<= 225 ;
          1800 : Address_next<= 450 ;
          1802 : Address_next<= 451 ;
          1803 : Address_next<= 225 ;
          1804 : Address_next<= 112 ;
          1806 : Address_next<= 113 ;
          1807 : Address_next<= 226 ;
          1808 : Address_next<= 452 ;
          1810 : Address_next<= 453 ;
          1811 : Address_next<= 226 ;
          1813 : Address_next<= 227 ;
          1814 : Address_next<= 454 ;
          1816 : Address_next<= 455 ;
          1817 : Address_next<= 227 ;
          1818 : Address_next<= 113 ;
          1819 : Address_next<= 56 ;
          1821 : Address_next<= 57 ;
          1822 : Address_next<= 114 ;
          1823 : Address_next<= 228 ;
          1824 : Address_next<= 456 ;
          1826 : Address_next<= 457 ;
          1827 : Address_next<= 228 ;
          1829 : Address_next<= 229 ;
          1830 : Address_next<= 458 ;
          1832 : Address_next<= 459 ;
          1833 : Address_next<= 229 ;
          1834 : Address_next<= 114 ;
          1836 : Address_next<= 115 ;
          1837 : Address_next<= 230 ;
          1838 : Address_next<= 460 ;
          1840 : Address_next<= 461 ;
          1841 : Address_next<= 230 ;
          1843 : Address_next<= 231 ;
          1844 : Address_next<= 462 ;
          1846 : Address_next<= 463 ;
          1847 : Address_next<= 231 ;
          1848 : Address_next<= 115 ;
          1849 : Address_next<= 57 ;
          1850 : Address_next<= 28 ;
          1852 : Address_next<= 29 ;
          1853 : Address_next<= 58 ;
          1854 : Address_next<= 116 ;
          1855 : Address_next<= 232 ;
          1856 : Address_next<= 464 ;
          1858 : Address_next<= 465 ;
          1859 : Address_next<= 232 ;
          1861 : Address_next<= 233 ;
          1862 : Address_next<= 466 ;
          1864 : Address_next<= 467 ;
          1865 : Address_next<= 233 ;
          1866 : Address_next<= 116 ;
          1868 : Address_next<= 117 ;
          1869 : Address_next<= 234 ;
          1870 : Address_next<= 468 ;
          1872 : Address_next<= 469 ;
          1873 : Address_next<= 234 ;
          1875 : Address_next<= 235 ;
          1876 : Address_next<= 470 ;
          1878 : Address_next<= 471 ;
          1879 : Address_next<= 235 ;
          1880 : Address_next<= 117 ;
          1881 : Address_next<= 58 ;
          1883 : Address_next<= 59 ;
          1884 : Address_next<= 118 ;
          1885 : Address_next<= 236 ;
          1886 : Address_next<= 472 ;
          1888 : Address_next<= 473 ;
          1889 : Address_next<= 236 ;
          1891 : Address_next<= 237 ;
          1892 : Address_next<= 474 ;
          1894 : Address_next<= 475 ;
          1895 : Address_next<= 237 ;
          1896 : Address_next<= 118 ;
          1898 : Address_next<= 119 ;
          1899 : Address_next<= 238 ;
          1900 : Address_next<= 476 ;
          1902 : Address_next<= 477 ;
          1903 : Address_next<= 238 ;
          1905 : Address_next<= 239 ;
          1906 : Address_next<= 478 ;
          1908 : Address_next<= 479 ;
          1909 : Address_next<= 239 ;
          1910 : Address_next<= 119 ;
          1911 : Address_next<= 59 ;
          1912 : Address_next<= 29 ;
          1913 : Address_next<= 14 ;
          1915 : Address_next<= 15 ;
          1916 : Address_next<= 30 ;
          1917 : Address_next<= 60 ;
          1918 : Address_next<= 120 ;
          1919 : Address_next<= 240 ;
          1920 : Address_next<= 480 ;
          1922 : Address_next<= 481 ;
          1923 : Address_next<= 240 ;
          1925 : Address_next<= 241 ;
          1926 : Address_next<= 482 ;
          1928 : Address_next<= 483 ;
          1929 : Address_next<= 241 ;
          1930 : Address_next<= 120 ;
          1932 : Address_next<= 121 ;
          1933 : Address_next<= 242 ;
          1934 : Address_next<= 484 ;
          1936 : Address_next<= 485 ;
          1937 : Address_next<= 242 ;
          1939 : Address_next<= 243 ;
          1940 : Address_next<= 486 ;
          1942 : Address_next<= 487 ;
          1943 : Address_next<= 243 ;
          1944 : Address_next<= 121 ;
          1945 : Address_next<= 60 ;
          1947 : Address_next<= 61 ;
          1948 : Address_next<= 122 ;
          1949 : Address_next<= 244 ;
          1950 : Address_next<= 488 ;
          1952 : Address_next<= 489 ;
          1953 : Address_next<= 244 ;
          1955 : Address_next<= 245 ;
          1956 : Address_next<= 490 ;
          1958 : Address_next<= 491 ;
          1959 : Address_next<= 245 ;
          1960 : Address_next<= 122 ;
          1962 : Address_next<= 123 ;
          1963 : Address_next<= 246 ;
          1964 : Address_next<= 492 ;
          1966 : Address_next<= 493 ;
          1967 : Address_next<= 246 ;
          1969 : Address_next<= 247 ;
          1970 : Address_next<= 494 ;
          1972 : Address_next<= 495 ;
          1973 : Address_next<= 247 ;
          1974 : Address_next<= 123 ;
          1975 : Address_next<= 61 ;
          1976 : Address_next<= 30 ;
          1978 : Address_next<= 31 ;
          1979 : Address_next<= 62 ;
          1980 : Address_next<= 124 ;
          1981 : Address_next<= 248 ;
          1982 : Address_next<= 496 ;
          1984 : Address_next<= 497 ;
          1985 : Address_next<= 248 ;
          1987 : Address_next<= 249 ;
          1988 : Address_next<= 498 ;
          1990 : Address_next<= 499 ;
          1991 : Address_next<= 249 ;
          1992 : Address_next<= 124 ;
          1994 : Address_next<= 125 ;
          1995 : Address_next<= 250 ;
          1996 : Address_next<= 500 ;
          1998 : Address_next<= 501 ;
          1999 : Address_next<= 250 ;
          2001 : Address_next<= 251 ;
          2002 : Address_next<= 502 ;
          2004 : Address_next<= 503 ;
          2005 : Address_next<= 251 ;
          2006 : Address_next<= 125 ;
          2007 : Address_next<= 62 ;
          2009 : Address_next<= 63 ;
          2010 : Address_next<= 126 ;
          2011 : Address_next<= 252 ;
          2012 : Address_next<= 504 ;
          2014 : Address_next<= 505 ;
          2015 : Address_next<= 252 ;
          2017 : Address_next<= 253 ;
          2018 : Address_next<= 506 ;
          2020 : Address_next<= 507 ;
          2021 : Address_next<= 253 ;
          2022 : Address_next<= 126 ;
          2024 : Address_next<= 127 ;
          2025 : Address_next<= 254 ;
          2026 : Address_next<= 508 ;
          2028 : Address_next<= 509 ;
          2029 : Address_next<= 254 ;
          2031 : Address_next<= 255 ;
          2032 : Address_next<= 510 ;
          2034 : Address_next<= 511 ;
          2035 : Address_next<= 255 ;
          2036 : Address_next<= 127 ;
          2037 : Address_next<= 63 ;
          2038 : Address_next<= 31 ;
          2039 : Address_next<= 15 ;
          2040 : Address_next<= 7 ;
          2041 : Address_next<= 3 ;
          2042 : Address_next<= 1 ;
       endcase
      end
      else begin
           L_Nv_next                     <=1024;
           L_opcode_next <= TYPE1;
           L_part_count_next <= 0;
           Address_next <= 0;
      end
end
end
endmodule


