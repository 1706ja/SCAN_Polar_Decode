module opcode #(parameter P = 128) (clk, rst, channel, I_program_counter,O_opcode, O_opcode_next, O_opcode_delay,
        O_Nv,O_Nv_next, O_part_count,O_part_count_next, O_address, O_address_next, O_opcode_before, O_Nv_before, O_bit_count);
        input clk,rst;
        input channel;
        input [15:0] I_program_counter;
        output [3:0] O_opcode,O_opcode_next, O_opcode_before, O_opcode_delay;
        output [10:0] O_Nv, O_Nv_next, O_Nv_before;
        output [3:0] O_part_count, O_part_count_next;
        output [9:0] O_address, O_address_next;
        output [12:0] O_bit_count;
        localparam TYPE1     = 4'b0000;
        localparam TYPE2     = 4'b0001;
        localparam BOTTOM    = 4'b0010;
        localparam TYPE3     = 4'b0011;
        localparam IDLE      = 4'b1011;

        reg [3:0] L_opcode, L_opcode_next, L_opcode_before, L_opcode_delay;
        reg [10:0] L_Nv,L_Nv_next,L_Nv_before, L_Nv_delay;
        reg [3:0] L_part_count, L_part_count_next, L_part_count_delay;
        reg [9:0] Address, Address_next, Address_delay;
        reg[12:0] L_bit_count;
        
        // assignment of outputs
        assign O_opcode = L_opcode;
        assign O_opcode_delay = L_opcode_delay;
        assign O_opcode_next = L_opcode_next;
        assign O_opcode_before = L_opcode_before;
        assign O_Nv = L_Nv;
        assign O_Nv_next = L_Nv_next;
        assign O_Nv_before = L_Nv_before;
        assign O_part_count = L_part_count;
        assign O_part_count_next = L_part_count_next;
        assign O_address = Address;
        assign O_address_next = Address_next;
        assign O_bit_count = L_bit_count;


        wire islast, oprand;
       assign islast = (L_Nv_next) > (2*P*(1+L_part_count_next));
       assign oprand = (L_opcode_next==TYPE1||L_opcode_next==TYPE2);

       always @(posedge clk)
     begin       
           if(!rst) begin
                L_Nv_before <= L_Nv;        
                L_Nv <= L_Nv_delay;
                L_Nv_delay <= L_Nv_next;

                L_opcode_before <= L_opcode;
                L_opcode <= L_opcode_delay;
                L_opcode_delay <= L_opcode_next;


                L_part_count <= L_part_count_delay;
                L_part_count_delay <= L_part_count_next;

//                Address_before <= Address;       
                L_bit_count <= (L_bit_count+2*(L_opcode==BOTTOM));

                Address <= Address_delay;
                Address_delay <= Address_next;
            end
            else begin
              L_bit_count <= 0;
              L_Nv                          <=1024; 
              L_Nv_before                          <=1024; 
              L_Nv_delay                          <=1024; 

              L_opcode_before <= TYPE1;
              L_opcode <= TYPE1;
              L_opcode_delay <= TYPE1;


              L_part_count <= 0;
              L_part_count_delay <= 0;

              Address <= 0;
              Address_delay <= 0;
            end
        end



        always @(posedge clk) begin
            if(rst) begin
            
            L_Nv_next                     <=1024;
            L_opcode_next <= TYPE1;
            L_part_count_next <= 0;
            // Address <= -1;
            Address_next <= 0;
            end
            else begin
           if (channel) begin
              case (L_Nv_next)
                1024 : L_Nv_next <= islast ? 1024 : 512;
                512 : L_Nv_next <= islast ?  512 : (oprand?256:1024);
                256 : L_Nv_next <= islast ? 256 : (oprand?128:512);
                128 : L_Nv_next <= oprand ? 64 : 256;
                64 : L_Nv_next <= oprand ? 32 : 128;
                32 : L_Nv_next <= oprand ? 16 : 64;
                16 : L_Nv_next <= oprand ? 8 : 32;
                8 : L_Nv_next <= oprand ? 4 : 16;
                4 : L_Nv_next <= oprand ? 2 : 8;
                2 : L_Nv_next <= 4;
                default: L_Nv_next <= 1024;
              endcase

              case (L_opcode_next)
                TYPE1 : L_opcode_next <= islast ? TYPE1 : ( (L_Nv_next==4) ? BOTTOM : TYPE1 );
                TYPE2 : L_opcode_next <= islast ? TYPE2 : ( (L_Nv_next==4) ? BOTTOM : TYPE1 );
                TYPE3 : L_opcode_next <= islast ? TYPE3 : ( (Address_next[0]) ? TYPE3 : TYPE2);
                BOTTOM : L_opcode_next <= Address_next[0] ? TYPE3 : TYPE2 ;
                default: L_opcode_next <= TYPE1;
              endcase

                case (L_part_count_next)
                  0 : L_part_count_next <= (L_Nv_next>2*P) ? 1 : 0;
                  1 : L_part_count_next <= (L_Nv_next>4*P) ? 2 : 0;
                  2 : L_part_count_next <= (L_Nv_next>4*P) ? 3 : 0;
                  3 : L_part_count_next <=  0;
                  // 4 : L_part_count_next <= (L_Nv_next>8*P) ? 5 : 0;
                  // 5 : L_part_count_next <= (L_Nv_next>8*P) ? 6 : 0;
                  // 6 : L_part_count_next <= (L_Nv_next>8*P) ? 7 : 0;
                  // 7 : L_part_count_next <= 0;
                  default: L_part_count_next <= 0;
                endcase


          


       case(I_program_counter)
          12 : Address_next<= 1 ;
          15 : Address_next<= 1 ;
          16 : Address_next<= 2 ;
          18 : Address_next<= 3 ;
          19 : Address_next<= 1 ;
          22 : Address_next<= 1 ;
          23 : Address_next<= 2 ;
          24 : Address_next<= 4 ;
          26 : Address_next<= 5 ;
          27 : Address_next<= 2 ;
          29 : Address_next<= 3 ;
          30 : Address_next<= 6 ;
          32 : Address_next<= 7 ;
          33 : Address_next<= 3 ;
          34 : Address_next<= 1 ;
          37 : Address_next<= 1 ;
          38 : Address_next<= 2 ;
          39 : Address_next<= 4 ;
          40 : Address_next<= 8 ;
          42 : Address_next<= 9 ;
          43 : Address_next<= 4 ;
          45 : Address_next<= 5 ;
          46 : Address_next<= 10 ;
          48 : Address_next<= 11 ;
          49 : Address_next<= 5 ;
          50 : Address_next<= 2 ;
          52 : Address_next<= 3 ;
          53 : Address_next<= 6 ;
          54 : Address_next<= 12 ;
          56 : Address_next<= 13 ;
          57 : Address_next<= 6 ;
          59 : Address_next<= 7 ;
          60 : Address_next<= 14 ;
          62 : Address_next<= 15 ;
          63 : Address_next<= 7 ;
          64 : Address_next<= 3 ;
          65 : Address_next<= 1 ;
          68 : Address_next<= 1 ;
          69 : Address_next<= 2 ;
          70 : Address_next<= 4 ;
          71 : Address_next<= 8 ;
          72 : Address_next<= 16 ;
          74 : Address_next<= 17 ;
          75 : Address_next<= 8 ;
          77 : Address_next<= 9 ;
          78 : Address_next<= 18 ;
          80 : Address_next<= 19 ;
          81 : Address_next<= 9 ;
          82 : Address_next<= 4 ;
          84 : Address_next<= 5 ;
          85 : Address_next<= 10 ;
          86 : Address_next<= 20 ;
          88 : Address_next<= 21 ;
          89 : Address_next<= 10 ;
          91 : Address_next<= 11 ;
          92 : Address_next<= 22 ;
          94 : Address_next<= 23 ;
          95 : Address_next<= 11 ;
          96 : Address_next<= 5 ;
          97 : Address_next<= 2 ;
          99 : Address_next<= 3 ;
          100 : Address_next<= 6 ;
          101 : Address_next<= 12 ;
          102 : Address_next<= 24 ;
          104 : Address_next<= 25 ;
          105 : Address_next<= 12 ;
          107 : Address_next<= 13 ;
          108 : Address_next<= 26 ;
          110 : Address_next<= 27 ;
          111 : Address_next<= 13 ;
          112 : Address_next<= 6 ;
          114 : Address_next<= 7 ;
          115 : Address_next<= 14 ;
          116 : Address_next<= 28 ;
          118 : Address_next<= 29 ;
          119 : Address_next<= 14 ;
          121 : Address_next<= 15 ;
          122 : Address_next<= 30 ;
          124 : Address_next<= 31 ;
          125 : Address_next<= 15 ;
          126 : Address_next<= 7 ;
          127 : Address_next<= 3 ;
          128 : Address_next<= 1 ;
          131 : Address_next<= 1 ;
          132 : Address_next<= 2 ;
          133 : Address_next<= 4 ;
          134 : Address_next<= 8 ;
          135 : Address_next<= 16 ;
          136 : Address_next<= 32 ;
          138 : Address_next<= 33 ;
          139 : Address_next<= 16 ;
          141 : Address_next<= 17 ;
          142 : Address_next<= 34 ;
          144 : Address_next<= 35 ;
          145 : Address_next<= 17 ;
          146 : Address_next<= 8 ;
          148 : Address_next<= 9 ;
          149 : Address_next<= 18 ;
          150 : Address_next<= 36 ;
          152 : Address_next<= 37 ;
          153 : Address_next<= 18 ;
          155 : Address_next<= 19 ;
          156 : Address_next<= 38 ;
          158 : Address_next<= 39 ;
          159 : Address_next<= 19 ;
          160 : Address_next<= 9 ;
          161 : Address_next<= 4 ;
          163 : Address_next<= 5 ;
          164 : Address_next<= 10 ;
          165 : Address_next<= 20 ;
          166 : Address_next<= 40 ;
          168 : Address_next<= 41 ;
          169 : Address_next<= 20 ;
          171 : Address_next<= 21 ;
          172 : Address_next<= 42 ;
          174 : Address_next<= 43 ;
          175 : Address_next<= 21 ;
          176 : Address_next<= 10 ;
          178 : Address_next<= 11 ;
          179 : Address_next<= 22 ;
          180 : Address_next<= 44 ;
          182 : Address_next<= 45 ;
          183 : Address_next<= 22 ;
          185 : Address_next<= 23 ;
          186 : Address_next<= 46 ;
          188 : Address_next<= 47 ;
          189 : Address_next<= 23 ;
          190 : Address_next<= 11 ;
          191 : Address_next<= 5 ;
          192 : Address_next<= 2 ;
          194 : Address_next<= 3 ;
          195 : Address_next<= 6 ;
          196 : Address_next<= 12 ;
          197 : Address_next<= 24 ;
          198 : Address_next<= 48 ;
          200 : Address_next<= 49 ;
          201 : Address_next<= 24 ;
          203 : Address_next<= 25 ;
          204 : Address_next<= 50 ;
          206 : Address_next<= 51 ;
          207 : Address_next<= 25 ;
          208 : Address_next<= 12 ;
          210 : Address_next<= 13 ;
          211 : Address_next<= 26 ;
          212 : Address_next<= 52 ;
          214 : Address_next<= 53 ;
          215 : Address_next<= 26 ;
          217 : Address_next<= 27 ;
          218 : Address_next<= 54 ;
          220 : Address_next<= 55 ;
          221 : Address_next<= 27 ;
          222 : Address_next<= 13 ;
          223 : Address_next<= 6 ;
          225 : Address_next<= 7 ;
          226 : Address_next<= 14 ;
          227 : Address_next<= 28 ;
          228 : Address_next<= 56 ;
          230 : Address_next<= 57 ;
          231 : Address_next<= 28 ;
          233 : Address_next<= 29 ;
          234 : Address_next<= 58 ;
          236 : Address_next<= 59 ;
          237 : Address_next<= 29 ;
          238 : Address_next<= 14 ;
          240 : Address_next<= 15 ;
          241 : Address_next<= 30 ;
          242 : Address_next<= 60 ;
          244 : Address_next<= 61 ;
          245 : Address_next<= 30 ;
          247 : Address_next<= 31 ;
          248 : Address_next<= 62 ;
          250 : Address_next<= 63 ;
          251 : Address_next<= 31 ;
          252 : Address_next<= 15 ;
          253 : Address_next<= 7 ;
          254 : Address_next<= 3 ;
          255 : Address_next<= 1 ;
          258 : Address_next<= 1 ;
          259 : Address_next<= 2 ;
          260 : Address_next<= 4 ;
          261 : Address_next<= 8 ;
          262 : Address_next<= 16 ;
          263 : Address_next<= 32 ;
          264 : Address_next<= 64 ;
          266 : Address_next<= 65 ;
          267 : Address_next<= 32 ;
          269 : Address_next<= 33 ;
          270 : Address_next<= 66 ;
          272 : Address_next<= 67 ;
          273 : Address_next<= 33 ;
          274 : Address_next<= 16 ;
          276 : Address_next<= 17 ;
          277 : Address_next<= 34 ;
          278 : Address_next<= 68 ;
          280 : Address_next<= 69 ;
          281 : Address_next<= 34 ;
          283 : Address_next<= 35 ;
          284 : Address_next<= 70 ;
          286 : Address_next<= 71 ;
          287 : Address_next<= 35 ;
          288 : Address_next<= 17 ;
          289 : Address_next<= 8 ;
          291 : Address_next<= 9 ;
          292 : Address_next<= 18 ;
          293 : Address_next<= 36 ;
          294 : Address_next<= 72 ;
          296 : Address_next<= 73 ;
          297 : Address_next<= 36 ;
          299 : Address_next<= 37 ;
          300 : Address_next<= 74 ;
          302 : Address_next<= 75 ;
          303 : Address_next<= 37 ;
          304 : Address_next<= 18 ;
          306 : Address_next<= 19 ;
          307 : Address_next<= 38 ;
          308 : Address_next<= 76 ;
          310 : Address_next<= 77 ;
          311 : Address_next<= 38 ;
          313 : Address_next<= 39 ;
          314 : Address_next<= 78 ;
          316 : Address_next<= 79 ;
          317 : Address_next<= 39 ;
          318 : Address_next<= 19 ;
          319 : Address_next<= 9 ;
          320 : Address_next<= 4 ;
          322 : Address_next<= 5 ;
          323 : Address_next<= 10 ;
          324 : Address_next<= 20 ;
          325 : Address_next<= 40 ;
          326 : Address_next<= 80 ;
          328 : Address_next<= 81 ;
          329 : Address_next<= 40 ;
          331 : Address_next<= 41 ;
          332 : Address_next<= 82 ;
          334 : Address_next<= 83 ;
          335 : Address_next<= 41 ;
          336 : Address_next<= 20 ;
          338 : Address_next<= 21 ;
          339 : Address_next<= 42 ;
          340 : Address_next<= 84 ;
          342 : Address_next<= 85 ;
          343 : Address_next<= 42 ;
          345 : Address_next<= 43 ;
          346 : Address_next<= 86 ;
          348 : Address_next<= 87 ;
          349 : Address_next<= 43 ;
          350 : Address_next<= 21 ;
          351 : Address_next<= 10 ;
          353 : Address_next<= 11 ;
          354 : Address_next<= 22 ;
          355 : Address_next<= 44 ;
          356 : Address_next<= 88 ;
          358 : Address_next<= 89 ;
          359 : Address_next<= 44 ;
          361 : Address_next<= 45 ;
          362 : Address_next<= 90 ;
          364 : Address_next<= 91 ;
          365 : Address_next<= 45 ;
          366 : Address_next<= 22 ;
          368 : Address_next<= 23 ;
          369 : Address_next<= 46 ;
          370 : Address_next<= 92 ;
          372 : Address_next<= 93 ;
          373 : Address_next<= 46 ;
          375 : Address_next<= 47 ;
          376 : Address_next<= 94 ;
          378 : Address_next<= 95 ;
          379 : Address_next<= 47 ;
          380 : Address_next<= 23 ;
          381 : Address_next<= 11 ;
          382 : Address_next<= 5 ;
          383 : Address_next<= 2 ;
          385 : Address_next<= 3 ;
          386 : Address_next<= 6 ;
          387 : Address_next<= 12 ;
          388 : Address_next<= 24 ;
          389 : Address_next<= 48 ;
          390 : Address_next<= 96 ;
          392 : Address_next<= 97 ;
          393 : Address_next<= 48 ;
          395 : Address_next<= 49 ;
          396 : Address_next<= 98 ;
          398 : Address_next<= 99 ;
          399 : Address_next<= 49 ;
          400 : Address_next<= 24 ;
          402 : Address_next<= 25 ;
          403 : Address_next<= 50 ;
          404 : Address_next<= 100 ;
          406 : Address_next<= 101 ;
          407 : Address_next<= 50 ;
          409 : Address_next<= 51 ;
          410 : Address_next<= 102 ;
          412 : Address_next<= 103 ;
          413 : Address_next<= 51 ;
          414 : Address_next<= 25 ;
          415 : Address_next<= 12 ;
          417 : Address_next<= 13 ;
          418 : Address_next<= 26 ;
          419 : Address_next<= 52 ;
          420 : Address_next<= 104 ;
          422 : Address_next<= 105 ;
          423 : Address_next<= 52 ;
          425 : Address_next<= 53 ;
          426 : Address_next<= 106 ;
          428 : Address_next<= 107 ;
          429 : Address_next<= 53 ;
          430 : Address_next<= 26 ;
          432 : Address_next<= 27 ;
          433 : Address_next<= 54 ;
          434 : Address_next<= 108 ;
          436 : Address_next<= 109 ;
          437 : Address_next<= 54 ;
          439 : Address_next<= 55 ;
          440 : Address_next<= 110 ;
          442 : Address_next<= 111 ;
          443 : Address_next<= 55 ;
          444 : Address_next<= 27 ;
          445 : Address_next<= 13 ;
          446 : Address_next<= 6 ;
          448 : Address_next<= 7 ;
          449 : Address_next<= 14 ;
          450 : Address_next<= 28 ;
          451 : Address_next<= 56 ;
          452 : Address_next<= 112 ;
          454 : Address_next<= 113 ;
          455 : Address_next<= 56 ;
          457 : Address_next<= 57 ;
          458 : Address_next<= 114 ;
          460 : Address_next<= 115 ;
          461 : Address_next<= 57 ;
          462 : Address_next<= 28 ;
          464 : Address_next<= 29 ;
          465 : Address_next<= 58 ;
          466 : Address_next<= 116 ;
          468 : Address_next<= 117 ;
          469 : Address_next<= 58 ;
          471 : Address_next<= 59 ;
          472 : Address_next<= 118 ;
          474 : Address_next<= 119 ;
          475 : Address_next<= 59 ;
          476 : Address_next<= 29 ;
          477 : Address_next<= 14 ;
          479 : Address_next<= 15 ;
          480 : Address_next<= 30 ;
          481 : Address_next<= 60 ;
          482 : Address_next<= 120 ;
          484 : Address_next<= 121 ;
          485 : Address_next<= 60 ;
          487 : Address_next<= 61 ;
          488 : Address_next<= 122 ;
          490 : Address_next<= 123 ;
          491 : Address_next<= 61 ;
          492 : Address_next<= 30 ;
          494 : Address_next<= 31 ;
          495 : Address_next<= 62 ;
          496 : Address_next<= 124 ;
          498 : Address_next<= 125 ;
          499 : Address_next<= 62 ;
          501 : Address_next<= 63 ;
          502 : Address_next<= 126 ;
          504 : Address_next<= 127 ;
          505 : Address_next<= 63 ;
          506 : Address_next<= 31 ;
          507 : Address_next<= 15 ;
          508 : Address_next<= 7 ;
          509 : Address_next<= 3 ;
          510 : Address_next<= 1 ;
          514 : Address_next<= 1 ;
          515 : Address_next<= 2 ;
          516 : Address_next<= 4 ;
          517 : Address_next<= 8 ;
          518 : Address_next<= 16 ;
          519 : Address_next<= 32 ;
          520 : Address_next<= 64 ;
          521 : Address_next<= 128 ;
          523 : Address_next<= 129 ;
          524 : Address_next<= 64 ;
          526 : Address_next<= 65 ;
          527 : Address_next<= 130 ;
          529 : Address_next<= 131 ;
          530 : Address_next<= 65 ;
          531 : Address_next<= 32 ;
          533 : Address_next<= 33 ;
          534 : Address_next<= 66 ;
          535 : Address_next<= 132 ;
          537 : Address_next<= 133 ;
          538 : Address_next<= 66 ;
          540 : Address_next<= 67 ;
          541 : Address_next<= 134 ;
          543 : Address_next<= 135 ;
          544 : Address_next<= 67 ;
          545 : Address_next<= 33 ;
          546 : Address_next<= 16 ;
          548 : Address_next<= 17 ;
          549 : Address_next<= 34 ;
          550 : Address_next<= 68 ;
          551 : Address_next<= 136 ;
          553 : Address_next<= 137 ;
          554 : Address_next<= 68 ;
          556 : Address_next<= 69 ;
          557 : Address_next<= 138 ;
          559 : Address_next<= 139 ;
          560 : Address_next<= 69 ;
          561 : Address_next<= 34 ;
          563 : Address_next<= 35 ;
          564 : Address_next<= 70 ;
          565 : Address_next<= 140 ;
          567 : Address_next<= 141 ;
          568 : Address_next<= 70 ;
          570 : Address_next<= 71 ;
          571 : Address_next<= 142 ;
          573 : Address_next<= 143 ;
          574 : Address_next<= 71 ;
          575 : Address_next<= 35 ;
          576 : Address_next<= 17 ;
          577 : Address_next<= 8 ;
          579 : Address_next<= 9 ;
          580 : Address_next<= 18 ;
          581 : Address_next<= 36 ;
          582 : Address_next<= 72 ;
          583 : Address_next<= 144 ;
          585 : Address_next<= 145 ;
          586 : Address_next<= 72 ;
          588 : Address_next<= 73 ;
          589 : Address_next<= 146 ;
          591 : Address_next<= 147 ;
          592 : Address_next<= 73 ;
          593 : Address_next<= 36 ;
          595 : Address_next<= 37 ;
          596 : Address_next<= 74 ;
          597 : Address_next<= 148 ;
          599 : Address_next<= 149 ;
          600 : Address_next<= 74 ;
          602 : Address_next<= 75 ;
          603 : Address_next<= 150 ;
          605 : Address_next<= 151 ;
          606 : Address_next<= 75 ;
          607 : Address_next<= 37 ;
          608 : Address_next<= 18 ;
          610 : Address_next<= 19 ;
          611 : Address_next<= 38 ;
          612 : Address_next<= 76 ;
          613 : Address_next<= 152 ;
          615 : Address_next<= 153 ;
          616 : Address_next<= 76 ;
          618 : Address_next<= 77 ;
          619 : Address_next<= 154 ;
          621 : Address_next<= 155 ;
          622 : Address_next<= 77 ;
          623 : Address_next<= 38 ;
          625 : Address_next<= 39 ;
          626 : Address_next<= 78 ;
          627 : Address_next<= 156 ;
          629 : Address_next<= 157 ;
          630 : Address_next<= 78 ;
          632 : Address_next<= 79 ;
          633 : Address_next<= 158 ;
          635 : Address_next<= 159 ;
          636 : Address_next<= 79 ;
          637 : Address_next<= 39 ;
          638 : Address_next<= 19 ;
          639 : Address_next<= 9 ;
          640 : Address_next<= 4 ;
          642 : Address_next<= 5 ;
          643 : Address_next<= 10 ;
          644 : Address_next<= 20 ;
          645 : Address_next<= 40 ;
          646 : Address_next<= 80 ;
          647 : Address_next<= 160 ;
          649 : Address_next<= 161 ;
          650 : Address_next<= 80 ;
          652 : Address_next<= 81 ;
          653 : Address_next<= 162 ;
          655 : Address_next<= 163 ;
          656 : Address_next<= 81 ;
          657 : Address_next<= 40 ;
          659 : Address_next<= 41 ;
          660 : Address_next<= 82 ;
          661 : Address_next<= 164 ;
          663 : Address_next<= 165 ;
          664 : Address_next<= 82 ;
          666 : Address_next<= 83 ;
          667 : Address_next<= 166 ;
          669 : Address_next<= 167 ;
          670 : Address_next<= 83 ;
          671 : Address_next<= 41 ;
          672 : Address_next<= 20 ;
          674 : Address_next<= 21 ;
          675 : Address_next<= 42 ;
          676 : Address_next<= 84 ;
          677 : Address_next<= 168 ;
          679 : Address_next<= 169 ;
          680 : Address_next<= 84 ;
          682 : Address_next<= 85 ;
          683 : Address_next<= 170 ;
          685 : Address_next<= 171 ;
          686 : Address_next<= 85 ;
          687 : Address_next<= 42 ;
          689 : Address_next<= 43 ;
          690 : Address_next<= 86 ;
          691 : Address_next<= 172 ;
          693 : Address_next<= 173 ;
          694 : Address_next<= 86 ;
          696 : Address_next<= 87 ;
          697 : Address_next<= 174 ;
          699 : Address_next<= 175 ;
          700 : Address_next<= 87 ;
          701 : Address_next<= 43 ;
          702 : Address_next<= 21 ;
          703 : Address_next<= 10 ;
          705 : Address_next<= 11 ;
          706 : Address_next<= 22 ;
          707 : Address_next<= 44 ;
          708 : Address_next<= 88 ;
          709 : Address_next<= 176 ;
          711 : Address_next<= 177 ;
          712 : Address_next<= 88 ;
          714 : Address_next<= 89 ;
          715 : Address_next<= 178 ;
          717 : Address_next<= 179 ;
          718 : Address_next<= 89 ;
          719 : Address_next<= 44 ;
          721 : Address_next<= 45 ;
          722 : Address_next<= 90 ;
          723 : Address_next<= 180 ;
          725 : Address_next<= 181 ;
          726 : Address_next<= 90 ;
          728 : Address_next<= 91 ;
          729 : Address_next<= 182 ;
          731 : Address_next<= 183 ;
          732 : Address_next<= 91 ;
          733 : Address_next<= 45 ;
          734 : Address_next<= 22 ;
          736 : Address_next<= 23 ;
          737 : Address_next<= 46 ;
          738 : Address_next<= 92 ;
          739 : Address_next<= 184 ;
          741 : Address_next<= 185 ;
          742 : Address_next<= 92 ;
          744 : Address_next<= 93 ;
          745 : Address_next<= 186 ;
          747 : Address_next<= 187 ;
          748 : Address_next<= 93 ;
          749 : Address_next<= 46 ;
          751 : Address_next<= 47 ;
          752 : Address_next<= 94 ;
          753 : Address_next<= 188 ;
          755 : Address_next<= 189 ;
          756 : Address_next<= 94 ;
          758 : Address_next<= 95 ;
          759 : Address_next<= 190 ;
          761 : Address_next<= 191 ;
          762 : Address_next<= 95 ;
          763 : Address_next<= 47 ;
          764 : Address_next<= 23 ;
          765 : Address_next<= 11 ;
          766 : Address_next<= 5 ;
          767 : Address_next<= 2 ;
          769 : Address_next<= 3 ;
          770 : Address_next<= 6 ;
          771 : Address_next<= 12 ;
          772 : Address_next<= 24 ;
          773 : Address_next<= 48 ;
          774 : Address_next<= 96 ;
          775 : Address_next<= 192 ;
          777 : Address_next<= 193 ;
          778 : Address_next<= 96 ;
          780 : Address_next<= 97 ;
          781 : Address_next<= 194 ;
          783 : Address_next<= 195 ;
          784 : Address_next<= 97 ;
          785 : Address_next<= 48 ;
          787 : Address_next<= 49 ;
          788 : Address_next<= 98 ;
          789 : Address_next<= 196 ;
          791 : Address_next<= 197 ;
          792 : Address_next<= 98 ;
          794 : Address_next<= 99 ;
          795 : Address_next<= 198 ;
          797 : Address_next<= 199 ;
          798 : Address_next<= 99 ;
          799 : Address_next<= 49 ;
          800 : Address_next<= 24 ;
          802 : Address_next<= 25 ;
          803 : Address_next<= 50 ;
          804 : Address_next<= 100 ;
          805 : Address_next<= 200 ;
          807 : Address_next<= 201 ;
          808 : Address_next<= 100 ;
          810 : Address_next<= 101 ;
          811 : Address_next<= 202 ;
          813 : Address_next<= 203 ;
          814 : Address_next<= 101 ;
          815 : Address_next<= 50 ;
          817 : Address_next<= 51 ;
          818 : Address_next<= 102 ;
          819 : Address_next<= 204 ;
          821 : Address_next<= 205 ;
          822 : Address_next<= 102 ;
          824 : Address_next<= 103 ;
          825 : Address_next<= 206 ;
          827 : Address_next<= 207 ;
          828 : Address_next<= 103 ;
          829 : Address_next<= 51 ;
          830 : Address_next<= 25 ;
          831 : Address_next<= 12 ;
          833 : Address_next<= 13 ;
          834 : Address_next<= 26 ;
          835 : Address_next<= 52 ;
          836 : Address_next<= 104 ;
          837 : Address_next<= 208 ;
          839 : Address_next<= 209 ;
          840 : Address_next<= 104 ;
          842 : Address_next<= 105 ;
          843 : Address_next<= 210 ;
          845 : Address_next<= 211 ;
          846 : Address_next<= 105 ;
          847 : Address_next<= 52 ;
          849 : Address_next<= 53 ;
          850 : Address_next<= 106 ;
          851 : Address_next<= 212 ;
          853 : Address_next<= 213 ;
          854 : Address_next<= 106 ;
          856 : Address_next<= 107 ;
          857 : Address_next<= 214 ;
          859 : Address_next<= 215 ;
          860 : Address_next<= 107 ;
          861 : Address_next<= 53 ;
          862 : Address_next<= 26 ;
          864 : Address_next<= 27 ;
          865 : Address_next<= 54 ;
          866 : Address_next<= 108 ;
          867 : Address_next<= 216 ;
          869 : Address_next<= 217 ;
          870 : Address_next<= 108 ;
          872 : Address_next<= 109 ;
          873 : Address_next<= 218 ;
          875 : Address_next<= 219 ;
          876 : Address_next<= 109 ;
          877 : Address_next<= 54 ;
          879 : Address_next<= 55 ;
          880 : Address_next<= 110 ;
          881 : Address_next<= 220 ;
          883 : Address_next<= 221 ;
          884 : Address_next<= 110 ;
          886 : Address_next<= 111 ;
          887 : Address_next<= 222 ;
          889 : Address_next<= 223 ;
          890 : Address_next<= 111 ;
          891 : Address_next<= 55 ;
          892 : Address_next<= 27 ;
          893 : Address_next<= 13 ;
          894 : Address_next<= 6 ;
          896 : Address_next<= 7 ;
          897 : Address_next<= 14 ;
          898 : Address_next<= 28 ;
          899 : Address_next<= 56 ;
          900 : Address_next<= 112 ;
          901 : Address_next<= 224 ;
          903 : Address_next<= 225 ;
          904 : Address_next<= 112 ;
          906 : Address_next<= 113 ;
          907 : Address_next<= 226 ;
          909 : Address_next<= 227 ;
          910 : Address_next<= 113 ;
          911 : Address_next<= 56 ;
          913 : Address_next<= 57 ;
          914 : Address_next<= 114 ;
          915 : Address_next<= 228 ;
          917 : Address_next<= 229 ;
          918 : Address_next<= 114 ;
          920 : Address_next<= 115 ;
          921 : Address_next<= 230 ;
          923 : Address_next<= 231 ;
          924 : Address_next<= 115 ;
          925 : Address_next<= 57 ;
          926 : Address_next<= 28 ;
          928 : Address_next<= 29 ;
          929 : Address_next<= 58 ;
          930 : Address_next<= 116 ;
          931 : Address_next<= 232 ;
          933 : Address_next<= 233 ;
          934 : Address_next<= 116 ;
          936 : Address_next<= 117 ;
          937 : Address_next<= 234 ;
          939 : Address_next<= 235 ;
          940 : Address_next<= 117 ;
          941 : Address_next<= 58 ;
          943 : Address_next<= 59 ;
          944 : Address_next<= 118 ;
          945 : Address_next<= 236 ;
          947 : Address_next<= 237 ;
          948 : Address_next<= 118 ;
          950 : Address_next<= 119 ;
          951 : Address_next<= 238 ;
          953 : Address_next<= 239 ;
          954 : Address_next<= 119 ;
          955 : Address_next<= 59 ;
          956 : Address_next<= 29 ;
          957 : Address_next<= 14 ;
          959 : Address_next<= 15 ;
          960 : Address_next<= 30 ;
          961 : Address_next<= 60 ;
          962 : Address_next<= 120 ;
          963 : Address_next<= 240 ;
          965 : Address_next<= 241 ;
          966 : Address_next<= 120 ;
          968 : Address_next<= 121 ;
          969 : Address_next<= 242 ;
          971 : Address_next<= 243 ;
          972 : Address_next<= 121 ;
          973 : Address_next<= 60 ;
          975 : Address_next<= 61 ;
          976 : Address_next<= 122 ;
          977 : Address_next<= 244 ;
          979 : Address_next<= 245 ;
          980 : Address_next<= 122 ;
          982 : Address_next<= 123 ;
          983 : Address_next<= 246 ;
          985 : Address_next<= 247 ;
          986 : Address_next<= 123 ;
          987 : Address_next<= 61 ;
          988 : Address_next<= 30 ;
          990 : Address_next<= 31 ;
          991 : Address_next<= 62 ;
          992 : Address_next<= 124 ;
          993 : Address_next<= 248 ;
          995 : Address_next<= 249 ;
          996 : Address_next<= 124 ;
          998 : Address_next<= 125 ;
          999 : Address_next<= 250 ;
          1001 : Address_next<= 251 ;
          1002 : Address_next<= 125 ;
          1003 : Address_next<= 62 ;
          1005 : Address_next<= 63 ;
          1006 : Address_next<= 126 ;
          1007 : Address_next<= 252 ;
          1009 : Address_next<= 253 ;
          1010 : Address_next<= 126 ;
          1012 : Address_next<= 127 ;
          1013 : Address_next<= 254 ;
          1015 : Address_next<= 255 ;
          1016 : Address_next<= 127 ;
          1017 : Address_next<= 63 ;
          1018 : Address_next<= 31 ;
          1019 : Address_next<= 15 ;
          1020 : Address_next<= 7 ;
          1021 : Address_next<= 3 ;
          1022 : Address_next<= 1 ;
          1029 : Address_next<= 1 ;
          1030 : Address_next<= 1 ;
          1031 : Address_next<= 2 ;
          1032 : Address_next<= 4 ;
          1033 : Address_next<= 8 ;
          1034 : Address_next<= 16 ;
          1035 : Address_next<= 32 ;
          1036 : Address_next<= 64 ;
          1037 : Address_next<= 128 ;
          1038 : Address_next<= 256 ;
          1040 : Address_next<= 257 ;
          1041 : Address_next<= 128 ;
          1043 : Address_next<= 129 ;
          1044 : Address_next<= 258 ;
          1046 : Address_next<= 259 ;
          1047 : Address_next<= 129 ;
          1048 : Address_next<= 64 ;
          1050 : Address_next<= 65 ;
          1051 : Address_next<= 130 ;
          1052 : Address_next<= 260 ;
          1054 : Address_next<= 261 ;
          1055 : Address_next<= 130 ;
          1057 : Address_next<= 131 ;
          1058 : Address_next<= 262 ;
          1060 : Address_next<= 263 ;
          1061 : Address_next<= 131 ;
          1062 : Address_next<= 65 ;
          1063 : Address_next<= 32 ;
          1065 : Address_next<= 33 ;
          1066 : Address_next<= 66 ;
          1067 : Address_next<= 132 ;
          1068 : Address_next<= 264 ;
          1070 : Address_next<= 265 ;
          1071 : Address_next<= 132 ;
          1073 : Address_next<= 133 ;
          1074 : Address_next<= 266 ;
          1076 : Address_next<= 267 ;
          1077 : Address_next<= 133 ;
          1078 : Address_next<= 66 ;
          1080 : Address_next<= 67 ;
          1081 : Address_next<= 134 ;
          1082 : Address_next<= 268 ;
          1084 : Address_next<= 269 ;
          1085 : Address_next<= 134 ;
          1087 : Address_next<= 135 ;
          1088 : Address_next<= 270 ;
          1090 : Address_next<= 271 ;
          1091 : Address_next<= 135 ;
          1092 : Address_next<= 67 ;
          1093 : Address_next<= 33 ;
          1094 : Address_next<= 16 ;
          1096 : Address_next<= 17 ;
          1097 : Address_next<= 34 ;
          1098 : Address_next<= 68 ;
          1099 : Address_next<= 136 ;
          1100 : Address_next<= 272 ;
          1102 : Address_next<= 273 ;
          1103 : Address_next<= 136 ;
          1105 : Address_next<= 137 ;
          1106 : Address_next<= 274 ;
          1108 : Address_next<= 275 ;
          1109 : Address_next<= 137 ;
          1110 : Address_next<= 68 ;
          1112 : Address_next<= 69 ;
          1113 : Address_next<= 138 ;
          1114 : Address_next<= 276 ;
          1116 : Address_next<= 277 ;
          1117 : Address_next<= 138 ;
          1119 : Address_next<= 139 ;
          1120 : Address_next<= 278 ;
          1122 : Address_next<= 279 ;
          1123 : Address_next<= 139 ;
          1124 : Address_next<= 69 ;
          1125 : Address_next<= 34 ;
          1127 : Address_next<= 35 ;
          1128 : Address_next<= 70 ;
          1129 : Address_next<= 140 ;
          1130 : Address_next<= 280 ;
          1132 : Address_next<= 281 ;
          1133 : Address_next<= 140 ;
          1135 : Address_next<= 141 ;
          1136 : Address_next<= 282 ;
          1138 : Address_next<= 283 ;
          1139 : Address_next<= 141 ;
          1140 : Address_next<= 70 ;
          1142 : Address_next<= 71 ;
          1143 : Address_next<= 142 ;
          1144 : Address_next<= 284 ;
          1146 : Address_next<= 285 ;
          1147 : Address_next<= 142 ;
          1149 : Address_next<= 143 ;
          1150 : Address_next<= 286 ;
          1152 : Address_next<= 287 ;
          1153 : Address_next<= 143 ;
          1154 : Address_next<= 71 ;
          1155 : Address_next<= 35 ;
          1156 : Address_next<= 17 ;
          1157 : Address_next<= 8 ;
          1159 : Address_next<= 9 ;
          1160 : Address_next<= 18 ;
          1161 : Address_next<= 36 ;
          1162 : Address_next<= 72 ;
          1163 : Address_next<= 144 ;
          1164 : Address_next<= 288 ;
          1166 : Address_next<= 289 ;
          1167 : Address_next<= 144 ;
          1169 : Address_next<= 145 ;
          1170 : Address_next<= 290 ;
          1172 : Address_next<= 291 ;
          1173 : Address_next<= 145 ;
          1174 : Address_next<= 72 ;
          1176 : Address_next<= 73 ;
          1177 : Address_next<= 146 ;
          1178 : Address_next<= 292 ;
          1180 : Address_next<= 293 ;
          1181 : Address_next<= 146 ;
          1183 : Address_next<= 147 ;
          1184 : Address_next<= 294 ;
          1186 : Address_next<= 295 ;
          1187 : Address_next<= 147 ;
          1188 : Address_next<= 73 ;
          1189 : Address_next<= 36 ;
          1191 : Address_next<= 37 ;
          1192 : Address_next<= 74 ;
          1193 : Address_next<= 148 ;
          1194 : Address_next<= 296 ;
          1196 : Address_next<= 297 ;
          1197 : Address_next<= 148 ;
          1199 : Address_next<= 149 ;
          1200 : Address_next<= 298 ;
          1202 : Address_next<= 299 ;
          1203 : Address_next<= 149 ;
          1204 : Address_next<= 74 ;
          1206 : Address_next<= 75 ;
          1207 : Address_next<= 150 ;
          1208 : Address_next<= 300 ;
          1210 : Address_next<= 301 ;
          1211 : Address_next<= 150 ;
          1213 : Address_next<= 151 ;
          1214 : Address_next<= 302 ;
          1216 : Address_next<= 303 ;
          1217 : Address_next<= 151 ;
          1218 : Address_next<= 75 ;
          1219 : Address_next<= 37 ;
          1220 : Address_next<= 18 ;
          1222 : Address_next<= 19 ;
          1223 : Address_next<= 38 ;
          1224 : Address_next<= 76 ;
          1225 : Address_next<= 152 ;
          1226 : Address_next<= 304 ;
          1228 : Address_next<= 305 ;
          1229 : Address_next<= 152 ;
          1231 : Address_next<= 153 ;
          1232 : Address_next<= 306 ;
          1234 : Address_next<= 307 ;
          1235 : Address_next<= 153 ;
          1236 : Address_next<= 76 ;
          1238 : Address_next<= 77 ;
          1239 : Address_next<= 154 ;
          1240 : Address_next<= 308 ;
          1242 : Address_next<= 309 ;
          1243 : Address_next<= 154 ;
          1245 : Address_next<= 155 ;
          1246 : Address_next<= 310 ;
          1248 : Address_next<= 311 ;
          1249 : Address_next<= 155 ;
          1250 : Address_next<= 77 ;
          1251 : Address_next<= 38 ;
          1253 : Address_next<= 39 ;
          1254 : Address_next<= 78 ;
          1255 : Address_next<= 156 ;
          1256 : Address_next<= 312 ;
          1258 : Address_next<= 313 ;
          1259 : Address_next<= 156 ;
          1261 : Address_next<= 157 ;
          1262 : Address_next<= 314 ;
          1264 : Address_next<= 315 ;
          1265 : Address_next<= 157 ;
          1266 : Address_next<= 78 ;
          1268 : Address_next<= 79 ;
          1269 : Address_next<= 158 ;
          1270 : Address_next<= 316 ;
          1272 : Address_next<= 317 ;
          1273 : Address_next<= 158 ;
          1275 : Address_next<= 159 ;
          1276 : Address_next<= 318 ;
          1278 : Address_next<= 319 ;
          1279 : Address_next<= 159 ;
          1280 : Address_next<= 79 ;
          1281 : Address_next<= 39 ;
          1282 : Address_next<= 19 ;
          1283 : Address_next<= 9 ;
          1284 : Address_next<= 4 ;
          1286 : Address_next<= 5 ;
          1287 : Address_next<= 10 ;
          1288 : Address_next<= 20 ;
          1289 : Address_next<= 40 ;
          1290 : Address_next<= 80 ;
          1291 : Address_next<= 160 ;
          1292 : Address_next<= 320 ;
          1294 : Address_next<= 321 ;
          1295 : Address_next<= 160 ;
          1297 : Address_next<= 161 ;
          1298 : Address_next<= 322 ;
          1300 : Address_next<= 323 ;
          1301 : Address_next<= 161 ;
          1302 : Address_next<= 80 ;
          1304 : Address_next<= 81 ;
          1305 : Address_next<= 162 ;
          1306 : Address_next<= 324 ;
          1308 : Address_next<= 325 ;
          1309 : Address_next<= 162 ;
          1311 : Address_next<= 163 ;
          1312 : Address_next<= 326 ;
          1314 : Address_next<= 327 ;
          1315 : Address_next<= 163 ;
          1316 : Address_next<= 81 ;
          1317 : Address_next<= 40 ;
          1319 : Address_next<= 41 ;
          1320 : Address_next<= 82 ;
          1321 : Address_next<= 164 ;
          1322 : Address_next<= 328 ;
          1324 : Address_next<= 329 ;
          1325 : Address_next<= 164 ;
          1327 : Address_next<= 165 ;
          1328 : Address_next<= 330 ;
          1330 : Address_next<= 331 ;
          1331 : Address_next<= 165 ;
          1332 : Address_next<= 82 ;
          1334 : Address_next<= 83 ;
          1335 : Address_next<= 166 ;
          1336 : Address_next<= 332 ;
          1338 : Address_next<= 333 ;
          1339 : Address_next<= 166 ;
          1341 : Address_next<= 167 ;
          1342 : Address_next<= 334 ;
          1344 : Address_next<= 335 ;
          1345 : Address_next<= 167 ;
          1346 : Address_next<= 83 ;
          1347 : Address_next<= 41 ;
          1348 : Address_next<= 20 ;
          1350 : Address_next<= 21 ;
          1351 : Address_next<= 42 ;
          1352 : Address_next<= 84 ;
          1353 : Address_next<= 168 ;
          1354 : Address_next<= 336 ;
          1356 : Address_next<= 337 ;
          1357 : Address_next<= 168 ;
          1359 : Address_next<= 169 ;
          1360 : Address_next<= 338 ;
          1362 : Address_next<= 339 ;
          1363 : Address_next<= 169 ;
          1364 : Address_next<= 84 ;
          1366 : Address_next<= 85 ;
          1367 : Address_next<= 170 ;
          1368 : Address_next<= 340 ;
          1370 : Address_next<= 341 ;
          1371 : Address_next<= 170 ;
          1373 : Address_next<= 171 ;
          1374 : Address_next<= 342 ;
          1376 : Address_next<= 343 ;
          1377 : Address_next<= 171 ;
          1378 : Address_next<= 85 ;
          1379 : Address_next<= 42 ;
          1381 : Address_next<= 43 ;
          1382 : Address_next<= 86 ;
          1383 : Address_next<= 172 ;
          1384 : Address_next<= 344 ;
          1386 : Address_next<= 345 ;
          1387 : Address_next<= 172 ;
          1389 : Address_next<= 173 ;
          1390 : Address_next<= 346 ;
          1392 : Address_next<= 347 ;
          1393 : Address_next<= 173 ;
          1394 : Address_next<= 86 ;
          1396 : Address_next<= 87 ;
          1397 : Address_next<= 174 ;
          1398 : Address_next<= 348 ;
          1400 : Address_next<= 349 ;
          1401 : Address_next<= 174 ;
          1403 : Address_next<= 175 ;
          1404 : Address_next<= 350 ;
          1406 : Address_next<= 351 ;
          1407 : Address_next<= 175 ;
          1408 : Address_next<= 87 ;
          1409 : Address_next<= 43 ;
          1410 : Address_next<= 21 ;
          1411 : Address_next<= 10 ;
          1413 : Address_next<= 11 ;
          1414 : Address_next<= 22 ;
          1415 : Address_next<= 44 ;
          1416 : Address_next<= 88 ;
          1417 : Address_next<= 176 ;
          1418 : Address_next<= 352 ;
          1420 : Address_next<= 353 ;
          1421 : Address_next<= 176 ;
          1423 : Address_next<= 177 ;
          1424 : Address_next<= 354 ;
          1426 : Address_next<= 355 ;
          1427 : Address_next<= 177 ;
          1428 : Address_next<= 88 ;
          1430 : Address_next<= 89 ;
          1431 : Address_next<= 178 ;
          1432 : Address_next<= 356 ;
          1434 : Address_next<= 357 ;
          1435 : Address_next<= 178 ;
          1437 : Address_next<= 179 ;
          1438 : Address_next<= 358 ;
          1440 : Address_next<= 359 ;
          1441 : Address_next<= 179 ;
          1442 : Address_next<= 89 ;
          1443 : Address_next<= 44 ;
          1445 : Address_next<= 45 ;
          1446 : Address_next<= 90 ;
          1447 : Address_next<= 180 ;
          1448 : Address_next<= 360 ;
          1450 : Address_next<= 361 ;
          1451 : Address_next<= 180 ;
          1453 : Address_next<= 181 ;
          1454 : Address_next<= 362 ;
          1456 : Address_next<= 363 ;
          1457 : Address_next<= 181 ;
          1458 : Address_next<= 90 ;
          1460 : Address_next<= 91 ;
          1461 : Address_next<= 182 ;
          1462 : Address_next<= 364 ;
          1464 : Address_next<= 365 ;
          1465 : Address_next<= 182 ;
          1467 : Address_next<= 183 ;
          1468 : Address_next<= 366 ;
          1470 : Address_next<= 367 ;
          1471 : Address_next<= 183 ;
          1472 : Address_next<= 91 ;
          1473 : Address_next<= 45 ;
          1474 : Address_next<= 22 ;
          1476 : Address_next<= 23 ;
          1477 : Address_next<= 46 ;
          1478 : Address_next<= 92 ;
          1479 : Address_next<= 184 ;
          1480 : Address_next<= 368 ;
          1482 : Address_next<= 369 ;
          1483 : Address_next<= 184 ;
          1485 : Address_next<= 185 ;
          1486 : Address_next<= 370 ;
          1488 : Address_next<= 371 ;
          1489 : Address_next<= 185 ;
          1490 : Address_next<= 92 ;
          1492 : Address_next<= 93 ;
          1493 : Address_next<= 186 ;
          1494 : Address_next<= 372 ;
          1496 : Address_next<= 373 ;
          1497 : Address_next<= 186 ;
          1499 : Address_next<= 187 ;
          1500 : Address_next<= 374 ;
          1502 : Address_next<= 375 ;
          1503 : Address_next<= 187 ;
          1504 : Address_next<= 93 ;
          1505 : Address_next<= 46 ;
          1507 : Address_next<= 47 ;
          1508 : Address_next<= 94 ;
          1509 : Address_next<= 188 ;
          1510 : Address_next<= 376 ;
          1512 : Address_next<= 377 ;
          1513 : Address_next<= 188 ;
          1515 : Address_next<= 189 ;
          1516 : Address_next<= 378 ;
          1518 : Address_next<= 379 ;
          1519 : Address_next<= 189 ;
          1520 : Address_next<= 94 ;
          1522 : Address_next<= 95 ;
          1523 : Address_next<= 190 ;
          1524 : Address_next<= 380 ;
          1526 : Address_next<= 381 ;
          1527 : Address_next<= 190 ;
          1529 : Address_next<= 191 ;
          1530 : Address_next<= 382 ;
          1532 : Address_next<= 383 ;
          1533 : Address_next<= 191 ;
          1534 : Address_next<= 95 ;
          1535 : Address_next<= 47 ;
          1536 : Address_next<= 23 ;
          1537 : Address_next<= 11 ;
          1538 : Address_next<= 5 ;
          1539 : Address_next<= 2 ;
          1542 : Address_next<= 3 ;
          1543 : Address_next<= 6 ;
          1544 : Address_next<= 12 ;
          1545 : Address_next<= 24 ;
          1546 : Address_next<= 48 ;
          1547 : Address_next<= 96 ;
          1548 : Address_next<= 192 ;
          1549 : Address_next<= 384 ;
          1551 : Address_next<= 385 ;
          1552 : Address_next<= 192 ;
          1554 : Address_next<= 193 ;
          1555 : Address_next<= 386 ;
          1557 : Address_next<= 387 ;
          1558 : Address_next<= 193 ;
          1559 : Address_next<= 96 ;
          1561 : Address_next<= 97 ;
          1562 : Address_next<= 194 ;
          1563 : Address_next<= 388 ;
          1565 : Address_next<= 389 ;
          1566 : Address_next<= 194 ;
          1568 : Address_next<= 195 ;
          1569 : Address_next<= 390 ;
          1571 : Address_next<= 391 ;
          1572 : Address_next<= 195 ;
          1573 : Address_next<= 97 ;
          1574 : Address_next<= 48 ;
          1576 : Address_next<= 49 ;
          1577 : Address_next<= 98 ;
          1578 : Address_next<= 196 ;
          1579 : Address_next<= 392 ;
          1581 : Address_next<= 393 ;
          1582 : Address_next<= 196 ;
          1584 : Address_next<= 197 ;
          1585 : Address_next<= 394 ;
          1587 : Address_next<= 395 ;
          1588 : Address_next<= 197 ;
          1589 : Address_next<= 98 ;
          1591 : Address_next<= 99 ;
          1592 : Address_next<= 198 ;
          1593 : Address_next<= 396 ;
          1595 : Address_next<= 397 ;
          1596 : Address_next<= 198 ;
          1598 : Address_next<= 199 ;
          1599 : Address_next<= 398 ;
          1601 : Address_next<= 399 ;
          1602 : Address_next<= 199 ;
          1603 : Address_next<= 99 ;
          1604 : Address_next<= 49 ;
          1605 : Address_next<= 24 ;
          1607 : Address_next<= 25 ;
          1608 : Address_next<= 50 ;
          1609 : Address_next<= 100 ;
          1610 : Address_next<= 200 ;
          1611 : Address_next<= 400 ;
          1613 : Address_next<= 401 ;
          1614 : Address_next<= 200 ;
          1616 : Address_next<= 201 ;
          1617 : Address_next<= 402 ;
          1619 : Address_next<= 403 ;
          1620 : Address_next<= 201 ;
          1621 : Address_next<= 100 ;
          1623 : Address_next<= 101 ;
          1624 : Address_next<= 202 ;
          1625 : Address_next<= 404 ;
          1627 : Address_next<= 405 ;
          1628 : Address_next<= 202 ;
          1630 : Address_next<= 203 ;
          1631 : Address_next<= 406 ;
          1633 : Address_next<= 407 ;
          1634 : Address_next<= 203 ;
          1635 : Address_next<= 101 ;
          1636 : Address_next<= 50 ;
          1638 : Address_next<= 51 ;
          1639 : Address_next<= 102 ;
          1640 : Address_next<= 204 ;
          1641 : Address_next<= 408 ;
          1643 : Address_next<= 409 ;
          1644 : Address_next<= 204 ;
          1646 : Address_next<= 205 ;
          1647 : Address_next<= 410 ;
          1649 : Address_next<= 411 ;
          1650 : Address_next<= 205 ;
          1651 : Address_next<= 102 ;
          1653 : Address_next<= 103 ;
          1654 : Address_next<= 206 ;
          1655 : Address_next<= 412 ;
          1657 : Address_next<= 413 ;
          1658 : Address_next<= 206 ;
          1660 : Address_next<= 207 ;
          1661 : Address_next<= 414 ;
          1663 : Address_next<= 415 ;
          1664 : Address_next<= 207 ;
          1665 : Address_next<= 103 ;
          1666 : Address_next<= 51 ;
          1667 : Address_next<= 25 ;
          1668 : Address_next<= 12 ;
          1670 : Address_next<= 13 ;
          1671 : Address_next<= 26 ;
          1672 : Address_next<= 52 ;
          1673 : Address_next<= 104 ;
          1674 : Address_next<= 208 ;
          1675 : Address_next<= 416 ;
          1677 : Address_next<= 417 ;
          1678 : Address_next<= 208 ;
          1680 : Address_next<= 209 ;
          1681 : Address_next<= 418 ;
          1683 : Address_next<= 419 ;
          1684 : Address_next<= 209 ;
          1685 : Address_next<= 104 ;
          1687 : Address_next<= 105 ;
          1688 : Address_next<= 210 ;
          1689 : Address_next<= 420 ;
          1691 : Address_next<= 421 ;
          1692 : Address_next<= 210 ;
          1694 : Address_next<= 211 ;
          1695 : Address_next<= 422 ;
          1697 : Address_next<= 423 ;
          1698 : Address_next<= 211 ;
          1699 : Address_next<= 105 ;
          1700 : Address_next<= 52 ;
          1702 : Address_next<= 53 ;
          1703 : Address_next<= 106 ;
          1704 : Address_next<= 212 ;
          1705 : Address_next<= 424 ;
          1707 : Address_next<= 425 ;
          1708 : Address_next<= 212 ;
          1710 : Address_next<= 213 ;
          1711 : Address_next<= 426 ;
          1713 : Address_next<= 427 ;
          1714 : Address_next<= 213 ;
          1715 : Address_next<= 106 ;
          1717 : Address_next<= 107 ;
          1718 : Address_next<= 214 ;
          1719 : Address_next<= 428 ;
          1721 : Address_next<= 429 ;
          1722 : Address_next<= 214 ;
          1724 : Address_next<= 215 ;
          1725 : Address_next<= 430 ;
          1727 : Address_next<= 431 ;
          1728 : Address_next<= 215 ;
          1729 : Address_next<= 107 ;
          1730 : Address_next<= 53 ;
          1731 : Address_next<= 26 ;
          1733 : Address_next<= 27 ;
          1734 : Address_next<= 54 ;
          1735 : Address_next<= 108 ;
          1736 : Address_next<= 216 ;
          1737 : Address_next<= 432 ;
          1739 : Address_next<= 433 ;
          1740 : Address_next<= 216 ;
          1742 : Address_next<= 217 ;
          1743 : Address_next<= 434 ;
          1745 : Address_next<= 435 ;
          1746 : Address_next<= 217 ;
          1747 : Address_next<= 108 ;
          1749 : Address_next<= 109 ;
          1750 : Address_next<= 218 ;
          1751 : Address_next<= 436 ;
          1753 : Address_next<= 437 ;
          1754 : Address_next<= 218 ;
          1756 : Address_next<= 219 ;
          1757 : Address_next<= 438 ;
          1759 : Address_next<= 439 ;
          1760 : Address_next<= 219 ;
          1761 : Address_next<= 109 ;
          1762 : Address_next<= 54 ;
          1764 : Address_next<= 55 ;
          1765 : Address_next<= 110 ;
          1766 : Address_next<= 220 ;
          1767 : Address_next<= 440 ;
          1769 : Address_next<= 441 ;
          1770 : Address_next<= 220 ;
          1772 : Address_next<= 221 ;
          1773 : Address_next<= 442 ;
          1775 : Address_next<= 443 ;
          1776 : Address_next<= 221 ;
          1777 : Address_next<= 110 ;
          1779 : Address_next<= 111 ;
          1780 : Address_next<= 222 ;
          1781 : Address_next<= 444 ;
          1783 : Address_next<= 445 ;
          1784 : Address_next<= 222 ;
          1786 : Address_next<= 223 ;
          1787 : Address_next<= 446 ;
          1789 : Address_next<= 447 ;
          1790 : Address_next<= 223 ;
          1791 : Address_next<= 111 ;
          1792 : Address_next<= 55 ;
          1793 : Address_next<= 27 ;
          1794 : Address_next<= 13 ;
          1795 : Address_next<= 6 ;
          1797 : Address_next<= 7 ;
          1798 : Address_next<= 14 ;
          1799 : Address_next<= 28 ;
          1800 : Address_next<= 56 ;
          1801 : Address_next<= 112 ;
          1802 : Address_next<= 224 ;
          1803 : Address_next<= 448 ;
          1805 : Address_next<= 449 ;
          1806 : Address_next<= 224 ;
          1808 : Address_next<= 225 ;
          1809 : Address_next<= 450 ;
          1811 : Address_next<= 451 ;
          1812 : Address_next<= 225 ;
          1813 : Address_next<= 112 ;
          1815 : Address_next<= 113 ;
          1816 : Address_next<= 226 ;
          1817 : Address_next<= 452 ;
          1819 : Address_next<= 453 ;
          1820 : Address_next<= 226 ;
          1822 : Address_next<= 227 ;
          1823 : Address_next<= 454 ;
          1825 : Address_next<= 455 ;
          1826 : Address_next<= 227 ;
          1827 : Address_next<= 113 ;
          1828 : Address_next<= 56 ;
          1830 : Address_next<= 57 ;
          1831 : Address_next<= 114 ;
          1832 : Address_next<= 228 ;
          1833 : Address_next<= 456 ;
          1835 : Address_next<= 457 ;
          1836 : Address_next<= 228 ;
          1838 : Address_next<= 229 ;
          1839 : Address_next<= 458 ;
          1841 : Address_next<= 459 ;
          1842 : Address_next<= 229 ;
          1843 : Address_next<= 114 ;
          1845 : Address_next<= 115 ;
          1846 : Address_next<= 230 ;
          1847 : Address_next<= 460 ;
          1849 : Address_next<= 461 ;
          1850 : Address_next<= 230 ;
          1852 : Address_next<= 231 ;
          1853 : Address_next<= 462 ;
          1855 : Address_next<= 463 ;
          1856 : Address_next<= 231 ;
          1857 : Address_next<= 115 ;
          1858 : Address_next<= 57 ;
          1859 : Address_next<= 28 ;
          1861 : Address_next<= 29 ;
          1862 : Address_next<= 58 ;
          1863 : Address_next<= 116 ;
          1864 : Address_next<= 232 ;
          1865 : Address_next<= 464 ;
          1867 : Address_next<= 465 ;
          1868 : Address_next<= 232 ;
          1870 : Address_next<= 233 ;
          1871 : Address_next<= 466 ;
          1873 : Address_next<= 467 ;
          1874 : Address_next<= 233 ;
          1875 : Address_next<= 116 ;
          1877 : Address_next<= 117 ;
          1878 : Address_next<= 234 ;
          1879 : Address_next<= 468 ;
          1881 : Address_next<= 469 ;
          1882 : Address_next<= 234 ;
          1884 : Address_next<= 235 ;
          1885 : Address_next<= 470 ;
          1887 : Address_next<= 471 ;
          1888 : Address_next<= 235 ;
          1889 : Address_next<= 117 ;
          1890 : Address_next<= 58 ;
          1892 : Address_next<= 59 ;
          1893 : Address_next<= 118 ;
          1894 : Address_next<= 236 ;
          1895 : Address_next<= 472 ;
          1897 : Address_next<= 473 ;
          1898 : Address_next<= 236 ;
          1900 : Address_next<= 237 ;
          1901 : Address_next<= 474 ;
          1903 : Address_next<= 475 ;
          1904 : Address_next<= 237 ;
          1905 : Address_next<= 118 ;
          1907 : Address_next<= 119 ;
          1908 : Address_next<= 238 ;
          1909 : Address_next<= 476 ;
          1911 : Address_next<= 477 ;
          1912 : Address_next<= 238 ;
          1914 : Address_next<= 239 ;
          1915 : Address_next<= 478 ;
          1917 : Address_next<= 479 ;
          1918 : Address_next<= 239 ;
          1919 : Address_next<= 119 ;
          1920 : Address_next<= 59 ;
          1921 : Address_next<= 29 ;
          1922 : Address_next<= 14 ;
          1924 : Address_next<= 15 ;
          1925 : Address_next<= 30 ;
          1926 : Address_next<= 60 ;
          1927 : Address_next<= 120 ;
          1928 : Address_next<= 240 ;
          1929 : Address_next<= 480 ;
          1931 : Address_next<= 481 ;
          1932 : Address_next<= 240 ;
          1934 : Address_next<= 241 ;
          1935 : Address_next<= 482 ;
          1937 : Address_next<= 483 ;
          1938 : Address_next<= 241 ;
          1939 : Address_next<= 120 ;
          1941 : Address_next<= 121 ;
          1942 : Address_next<= 242 ;
          1943 : Address_next<= 484 ;
          1945 : Address_next<= 485 ;
          1946 : Address_next<= 242 ;
          1948 : Address_next<= 243 ;
          1949 : Address_next<= 486 ;
          1951 : Address_next<= 487 ;
          1952 : Address_next<= 243 ;
          1953 : Address_next<= 121 ;
          1954 : Address_next<= 60 ;
          1956 : Address_next<= 61 ;
          1957 : Address_next<= 122 ;
          1958 : Address_next<= 244 ;
          1959 : Address_next<= 488 ;
          1961 : Address_next<= 489 ;
          1962 : Address_next<= 244 ;
          1964 : Address_next<= 245 ;
          1965 : Address_next<= 490 ;
          1967 : Address_next<= 491 ;
          1968 : Address_next<= 245 ;
          1969 : Address_next<= 122 ;
          1971 : Address_next<= 123 ;
          1972 : Address_next<= 246 ;
          1973 : Address_next<= 492 ;
          1975 : Address_next<= 493 ;
          1976 : Address_next<= 246 ;
          1978 : Address_next<= 247 ;
          1979 : Address_next<= 494 ;
          1981 : Address_next<= 495 ;
          1982 : Address_next<= 247 ;
          1983 : Address_next<= 123 ;
          1984 : Address_next<= 61 ;
          1985 : Address_next<= 30 ;
          1987 : Address_next<= 31 ;
          1988 : Address_next<= 62 ;
          1989 : Address_next<= 124 ;
          1990 : Address_next<= 248 ;
          1991 : Address_next<= 496 ;
          1993 : Address_next<= 497 ;
          1994 : Address_next<= 248 ;
          1996 : Address_next<= 249 ;
          1997 : Address_next<= 498 ;
          1999 : Address_next<= 499 ;
          2000 : Address_next<= 249 ;
          2001 : Address_next<= 124 ;
          2003 : Address_next<= 125 ;
          2004 : Address_next<= 250 ;
          2005 : Address_next<= 500 ;
          2007 : Address_next<= 501 ;
          2008 : Address_next<= 250 ;
          2010 : Address_next<= 251 ;
          2011 : Address_next<= 502 ;
          2013 : Address_next<= 503 ;
          2014 : Address_next<= 251 ;
          2015 : Address_next<= 125 ;
          2016 : Address_next<= 62 ;
          2018 : Address_next<= 63 ;
          2019 : Address_next<= 126 ;
          2020 : Address_next<= 252 ;
          2021 : Address_next<= 504 ;
          2023 : Address_next<= 505 ;
          2024 : Address_next<= 252 ;
          2026 : Address_next<= 253 ;
          2027 : Address_next<= 506 ;
          2029 : Address_next<= 507 ;
          2030 : Address_next<= 253 ;
          2031 : Address_next<= 126 ;
          2033 : Address_next<= 127 ;
          2034 : Address_next<= 254 ;
          2035 : Address_next<= 508 ;
          2037 : Address_next<= 509 ;
          2038 : Address_next<= 254 ;
          2040 : Address_next<= 255 ;
          2041 : Address_next<= 510 ;
          2043 : Address_next<= 511 ;
          2044 : Address_next<= 255 ;
          2045 : Address_next<= 127 ;
          2046 : Address_next<= 63 ;
          2047 : Address_next<= 31 ;
          2048 : Address_next<= 15 ;
          2049 : Address_next<= 7 ;
          2050 : Address_next<= 3 ;
          2051 : Address_next<= 1 ;
          2052 : Address_next<= 1 ;
        default : Address_next <= 0;
       endcase








      end
      else begin
           L_Nv_next                     <=1024;
           L_opcode_next <= TYPE1;
           L_part_count_next <= 0;
           Address_next <= 0;
      end
end
end
endmodule


