module opcode #(parameter P = 64) (clk, rst, channel, I_program_counter,O_opcode, O_opcode_next, O_opcode_delay,
        O_Nv,O_Nv_next, O_part_count,O_part_count_next, O_address, O_address_next, O_opcode_before, O_Nv_before, O_bit_count);
        input clk,rst;
        input channel;
        input [15:0] I_program_counter;
        output [3:0] O_opcode,O_opcode_next, O_opcode_before, O_opcode_delay;
        output [10:0] O_Nv, O_Nv_next, O_Nv_before;
        output [3:0] O_part_count, O_part_count_next;
        output [9:0] O_address, O_address_next;
        output [12:0] O_bit_count;
        localparam TYPE1     = 4'b0000;
        localparam TYPE2     = 4'b0001;
        localparam BOTTOM    = 4'b0010;
        localparam TYPE3     = 4'b0011;
        localparam IDLE      = 4'b1011;

        reg [3:0] L_opcode, L_opcode_next, L_opcode_before, L_opcode_delay;
        reg [10:0] L_Nv,L_Nv_next,L_Nv_before, L_Nv_delay;
        reg [3:0] L_part_count, L_part_count_next, L_part_count_delay;
        reg [9:0] Address, Address_next, Address_delay;
        reg[12:0] L_bit_count;
        
        // assignment of outputs
        assign O_opcode = L_opcode;
        assign O_opcode_delay = L_opcode_delay;
        assign O_opcode_next = L_opcode_next;
        assign O_opcode_before = L_opcode_before;
        assign O_Nv = L_Nv;
        assign O_Nv_next = L_Nv_next;
        assign O_Nv_before = L_Nv_before;
        assign O_part_count = L_part_count;
        assign O_part_count_next = L_part_count_next;
        assign O_address = Address;
        assign O_address_next = Address_next;
        assign O_bit_count = L_bit_count;


        wire islast, oprand;
       assign islast = (L_Nv_next) > (2*P*(1+L_part_count_next));
       assign oprand = (L_opcode_next==TYPE1||L_opcode_next==TYPE2);

       always @(posedge clk)
     begin       
           if(!rst) begin
                L_Nv_before <= L_Nv;        
                L_Nv <= L_Nv_delay;
                L_Nv_delay <= L_Nv_next;

                L_opcode_before <= L_opcode;
                L_opcode <= L_opcode_delay;
                L_opcode_delay <= L_opcode_next;


                L_part_count <= L_part_count_delay;
                L_part_count_delay <= L_part_count_next;

//                Address_before <= Address;       
                L_bit_count <= (L_bit_count+2*(L_opcode==BOTTOM));

                Address <= Address_delay;
                Address_delay <= Address_next;
            end
            else begin
              L_bit_count <= 0;
              L_Nv                          <=1024; 
              L_Nv_before                          <=1024; 
              L_Nv_delay                          <=1024; 

              L_opcode_before <= TYPE1;
              L_opcode <= TYPE1;
              L_opcode_delay <= TYPE1;


              L_part_count <= 0;
              L_part_count_delay <= 0;

              Address <= 0;
              Address_delay <= 0;
            end
        end



        always @(posedge clk) begin
            if(rst) begin
            
            L_Nv_next                     <=1024;
            L_opcode_next <= TYPE1;
            L_part_count_next <= 0;
            // Address <= -1;
            Address_next <= 0;
            end
            else begin
           if (channel) begin
              case (L_Nv_next)
                1024 : L_Nv_next <= islast ? 1024 : 512;
                512 : L_Nv_next <= islast ?  512 : (oprand?256:1024);
                256 : L_Nv_next <= islast ? 256 : (oprand?128:512);
                128 : L_Nv_next <= oprand ? 64 : 256;
                64 : L_Nv_next <= oprand ? 32 : 128;
                32 : L_Nv_next <= oprand ? 16 : 64;
                16 : L_Nv_next <= oprand ? 8 : 32;
                8 : L_Nv_next <= oprand ? 4 : 16;
                4 : L_Nv_next <= oprand ? 2 : 8;
                2 : L_Nv_next <= 4;
                default: L_Nv_next <= 1024;
              endcase

              case (L_opcode_next)
                TYPE1 : L_opcode_next <= islast ? TYPE1 : ( (L_Nv_next==4) ? BOTTOM : TYPE1 );
                TYPE2 : L_opcode_next <= islast ? TYPE2 : ( (L_Nv_next==4) ? BOTTOM : TYPE1 );
                TYPE3 : begin
                  L_opcode_next <= islast ? TYPE3 : ( 
                     (L_Nv_next==512): TYPE1 :
                    ((Address_next[0]) ? TYPE3 : TYPE2)
                    );
                end
                 
                BOTTOM : L_opcode_next <= Address_next[0] ? TYPE3 : TYPE2 ;
                default: L_opcode_next <= TYPE1;
              endcase

              L_part_count_next <= islast ? L_part_count_next+1 : 0;

          



       case(I_program_counter)
          19 : Address_next<= 1 ;
          22 : Address_next<= 1 ;
          23 : Address_next<= 2 ;
          25 : Address_next<= 3 ;
          26 : Address_next<= 1 ;
          29 : Address_next<= 1 ;
          30 : Address_next<= 2 ;
          31 : Address_next<= 4 ;
          33 : Address_next<= 5 ;
          34 : Address_next<= 2 ;
          36 : Address_next<= 3 ;
          37 : Address_next<= 6 ;
          39 : Address_next<= 7 ;
          40 : Address_next<= 3 ;
          41 : Address_next<= 1 ;
          44 : Address_next<= 1 ;
          45 : Address_next<= 2 ;
          46 : Address_next<= 4 ;
          47 : Address_next<= 8 ;
          49 : Address_next<= 9 ;
          50 : Address_next<= 4 ;
          52 : Address_next<= 5 ;
          53 : Address_next<= 10 ;
          55 : Address_next<= 11 ;
          56 : Address_next<= 5 ;
          57 : Address_next<= 2 ;
          59 : Address_next<= 3 ;
          60 : Address_next<= 6 ;
          61 : Address_next<= 12 ;
          63 : Address_next<= 13 ;
          64 : Address_next<= 6 ;
          66 : Address_next<= 7 ;
          67 : Address_next<= 14 ;
          69 : Address_next<= 15 ;
          70 : Address_next<= 7 ;
          71 : Address_next<= 3 ;
          72 : Address_next<= 1 ;
          75 : Address_next<= 1 ;
          76 : Address_next<= 2 ;
          77 : Address_next<= 4 ;
          78 : Address_next<= 8 ;
          79 : Address_next<= 16 ;
          81 : Address_next<= 17 ;
          82 : Address_next<= 8 ;
          84 : Address_next<= 9 ;
          85 : Address_next<= 18 ;
          87 : Address_next<= 19 ;
          88 : Address_next<= 9 ;
          89 : Address_next<= 4 ;
          91 : Address_next<= 5 ;
          92 : Address_next<= 10 ;
          93 : Address_next<= 20 ;
          95 : Address_next<= 21 ;
          96 : Address_next<= 10 ;
          98 : Address_next<= 11 ;
          99 : Address_next<= 22 ;
          101 : Address_next<= 23 ;
          102 : Address_next<= 11 ;
          103 : Address_next<= 5 ;
          104 : Address_next<= 2 ;
          106 : Address_next<= 3 ;
          107 : Address_next<= 6 ;
          108 : Address_next<= 12 ;
          109 : Address_next<= 24 ;
          111 : Address_next<= 25 ;
          112 : Address_next<= 12 ;
          114 : Address_next<= 13 ;
          115 : Address_next<= 26 ;
          117 : Address_next<= 27 ;
          118 : Address_next<= 13 ;
          119 : Address_next<= 6 ;
          121 : Address_next<= 7 ;
          122 : Address_next<= 14 ;
          123 : Address_next<= 28 ;
          125 : Address_next<= 29 ;
          126 : Address_next<= 14 ;
          128 : Address_next<= 15 ;
          129 : Address_next<= 30 ;
          131 : Address_next<= 31 ;
          132 : Address_next<= 15 ;
          133 : Address_next<= 7 ;
          134 : Address_next<= 3 ;
          135 : Address_next<= 1 ;
          138 : Address_next<= 1 ;
          139 : Address_next<= 2 ;
          140 : Address_next<= 4 ;
          141 : Address_next<= 8 ;
          142 : Address_next<= 16 ;
          143 : Address_next<= 32 ;
          145 : Address_next<= 33 ;
          146 : Address_next<= 16 ;
          148 : Address_next<= 17 ;
          149 : Address_next<= 34 ;
          151 : Address_next<= 35 ;
          152 : Address_next<= 17 ;
          153 : Address_next<= 8 ;
          155 : Address_next<= 9 ;
          156 : Address_next<= 18 ;
          157 : Address_next<= 36 ;
          159 : Address_next<= 37 ;
          160 : Address_next<= 18 ;
          162 : Address_next<= 19 ;
          163 : Address_next<= 38 ;
          165 : Address_next<= 39 ;
          166 : Address_next<= 19 ;
          167 : Address_next<= 9 ;
          168 : Address_next<= 4 ;
          170 : Address_next<= 5 ;
          171 : Address_next<= 10 ;
          172 : Address_next<= 20 ;
          173 : Address_next<= 40 ;
          175 : Address_next<= 41 ;
          176 : Address_next<= 20 ;
          178 : Address_next<= 21 ;
          179 : Address_next<= 42 ;
          181 : Address_next<= 43 ;
          182 : Address_next<= 21 ;
          183 : Address_next<= 10 ;
          185 : Address_next<= 11 ;
          186 : Address_next<= 22 ;
          187 : Address_next<= 44 ;
          189 : Address_next<= 45 ;
          190 : Address_next<= 22 ;
          192 : Address_next<= 23 ;
          193 : Address_next<= 46 ;
          195 : Address_next<= 47 ;
          196 : Address_next<= 23 ;
          197 : Address_next<= 11 ;
          198 : Address_next<= 5 ;
          199 : Address_next<= 2 ;
          201 : Address_next<= 3 ;
          202 : Address_next<= 6 ;
          203 : Address_next<= 12 ;
          204 : Address_next<= 24 ;
          205 : Address_next<= 48 ;
          207 : Address_next<= 49 ;
          208 : Address_next<= 24 ;
          210 : Address_next<= 25 ;
          211 : Address_next<= 50 ;
          213 : Address_next<= 51 ;
          214 : Address_next<= 25 ;
          215 : Address_next<= 12 ;
          217 : Address_next<= 13 ;
          218 : Address_next<= 26 ;
          219 : Address_next<= 52 ;
          221 : Address_next<= 53 ;
          222 : Address_next<= 26 ;
          224 : Address_next<= 27 ;
          225 : Address_next<= 54 ;
          227 : Address_next<= 55 ;
          228 : Address_next<= 27 ;
          229 : Address_next<= 13 ;
          230 : Address_next<= 6 ;
          232 : Address_next<= 7 ;
          233 : Address_next<= 14 ;
          234 : Address_next<= 28 ;
          235 : Address_next<= 56 ;
          237 : Address_next<= 57 ;
          238 : Address_next<= 28 ;
          240 : Address_next<= 29 ;
          241 : Address_next<= 58 ;
          243 : Address_next<= 59 ;
          244 : Address_next<= 29 ;
          245 : Address_next<= 14 ;
          247 : Address_next<= 15 ;
          248 : Address_next<= 30 ;
          249 : Address_next<= 60 ;
          251 : Address_next<= 61 ;
          252 : Address_next<= 30 ;
          254 : Address_next<= 31 ;
          255 : Address_next<= 62 ;
          257 : Address_next<= 63 ;
          258 : Address_next<= 31 ;
          259 : Address_next<= 15 ;
          260 : Address_next<= 7 ;
          261 : Address_next<= 3 ;
          262 : Address_next<= 1 ;
          266 : Address_next<= 1 ;
          267 : Address_next<= 2 ;
          268 : Address_next<= 4 ;
          269 : Address_next<= 8 ;
          270 : Address_next<= 16 ;
          271 : Address_next<= 32 ;
          272 : Address_next<= 64 ;
          274 : Address_next<= 65 ;
          275 : Address_next<= 32 ;
          277 : Address_next<= 33 ;
          278 : Address_next<= 66 ;
          280 : Address_next<= 67 ;
          281 : Address_next<= 33 ;
          282 : Address_next<= 16 ;
          284 : Address_next<= 17 ;
          285 : Address_next<= 34 ;
          286 : Address_next<= 68 ;
          288 : Address_next<= 69 ;
          289 : Address_next<= 34 ;
          291 : Address_next<= 35 ;
          292 : Address_next<= 70 ;
          294 : Address_next<= 71 ;
          295 : Address_next<= 35 ;
          296 : Address_next<= 17 ;
          297 : Address_next<= 8 ;
          299 : Address_next<= 9 ;
          300 : Address_next<= 18 ;
          301 : Address_next<= 36 ;
          302 : Address_next<= 72 ;
          304 : Address_next<= 73 ;
          305 : Address_next<= 36 ;
          307 : Address_next<= 37 ;
          308 : Address_next<= 74 ;
          310 : Address_next<= 75 ;
          311 : Address_next<= 37 ;
          312 : Address_next<= 18 ;
          314 : Address_next<= 19 ;
          315 : Address_next<= 38 ;
          316 : Address_next<= 76 ;
          318 : Address_next<= 77 ;
          319 : Address_next<= 38 ;
          321 : Address_next<= 39 ;
          322 : Address_next<= 78 ;
          324 : Address_next<= 79 ;
          325 : Address_next<= 39 ;
          326 : Address_next<= 19 ;
          327 : Address_next<= 9 ;
          328 : Address_next<= 4 ;
          330 : Address_next<= 5 ;
          331 : Address_next<= 10 ;
          332 : Address_next<= 20 ;
          333 : Address_next<= 40 ;
          334 : Address_next<= 80 ;
          336 : Address_next<= 81 ;
          337 : Address_next<= 40 ;
          339 : Address_next<= 41 ;
          340 : Address_next<= 82 ;
          342 : Address_next<= 83 ;
          343 : Address_next<= 41 ;
          344 : Address_next<= 20 ;
          346 : Address_next<= 21 ;
          347 : Address_next<= 42 ;
          348 : Address_next<= 84 ;
          350 : Address_next<= 85 ;
          351 : Address_next<= 42 ;
          353 : Address_next<= 43 ;
          354 : Address_next<= 86 ;
          356 : Address_next<= 87 ;
          357 : Address_next<= 43 ;
          358 : Address_next<= 21 ;
          359 : Address_next<= 10 ;
          361 : Address_next<= 11 ;
          362 : Address_next<= 22 ;
          363 : Address_next<= 44 ;
          364 : Address_next<= 88 ;
          366 : Address_next<= 89 ;
          367 : Address_next<= 44 ;
          369 : Address_next<= 45 ;
          370 : Address_next<= 90 ;
          372 : Address_next<= 91 ;
          373 : Address_next<= 45 ;
          374 : Address_next<= 22 ;
          376 : Address_next<= 23 ;
          377 : Address_next<= 46 ;
          378 : Address_next<= 92 ;
          380 : Address_next<= 93 ;
          381 : Address_next<= 46 ;
          383 : Address_next<= 47 ;
          384 : Address_next<= 94 ;
          386 : Address_next<= 95 ;
          387 : Address_next<= 47 ;
          388 : Address_next<= 23 ;
          389 : Address_next<= 11 ;
          390 : Address_next<= 5 ;
          391 : Address_next<= 2 ;
          393 : Address_next<= 3 ;
          394 : Address_next<= 6 ;
          395 : Address_next<= 12 ;
          396 : Address_next<= 24 ;
          397 : Address_next<= 48 ;
          398 : Address_next<= 96 ;
          400 : Address_next<= 97 ;
          401 : Address_next<= 48 ;
          403 : Address_next<= 49 ;
          404 : Address_next<= 98 ;
          406 : Address_next<= 99 ;
          407 : Address_next<= 49 ;
          408 : Address_next<= 24 ;
          410 : Address_next<= 25 ;
          411 : Address_next<= 50 ;
          412 : Address_next<= 100 ;
          414 : Address_next<= 101 ;
          415 : Address_next<= 50 ;
          417 : Address_next<= 51 ;
          418 : Address_next<= 102 ;
          420 : Address_next<= 103 ;
          421 : Address_next<= 51 ;
          422 : Address_next<= 25 ;
          423 : Address_next<= 12 ;
          425 : Address_next<= 13 ;
          426 : Address_next<= 26 ;
          427 : Address_next<= 52 ;
          428 : Address_next<= 104 ;
          430 : Address_next<= 105 ;
          431 : Address_next<= 52 ;
          433 : Address_next<= 53 ;
          434 : Address_next<= 106 ;
          436 : Address_next<= 107 ;
          437 : Address_next<= 53 ;
          438 : Address_next<= 26 ;
          440 : Address_next<= 27 ;
          441 : Address_next<= 54 ;
          442 : Address_next<= 108 ;
          444 : Address_next<= 109 ;
          445 : Address_next<= 54 ;
          447 : Address_next<= 55 ;
          448 : Address_next<= 110 ;
          450 : Address_next<= 111 ;
          451 : Address_next<= 55 ;
          452 : Address_next<= 27 ;
          453 : Address_next<= 13 ;
          454 : Address_next<= 6 ;
          456 : Address_next<= 7 ;
          457 : Address_next<= 14 ;
          458 : Address_next<= 28 ;
          459 : Address_next<= 56 ;
          460 : Address_next<= 112 ;
          462 : Address_next<= 113 ;
          463 : Address_next<= 56 ;
          465 : Address_next<= 57 ;
          466 : Address_next<= 114 ;
          468 : Address_next<= 115 ;
          469 : Address_next<= 57 ;
          470 : Address_next<= 28 ;
          472 : Address_next<= 29 ;
          473 : Address_next<= 58 ;
          474 : Address_next<= 116 ;
          476 : Address_next<= 117 ;
          477 : Address_next<= 58 ;
          479 : Address_next<= 59 ;
          480 : Address_next<= 118 ;
          482 : Address_next<= 119 ;
          483 : Address_next<= 59 ;
          484 : Address_next<= 29 ;
          485 : Address_next<= 14 ;
          487 : Address_next<= 15 ;
          488 : Address_next<= 30 ;
          489 : Address_next<= 60 ;
          490 : Address_next<= 120 ;
          492 : Address_next<= 121 ;
          493 : Address_next<= 60 ;
          495 : Address_next<= 61 ;
          496 : Address_next<= 122 ;
          498 : Address_next<= 123 ;
          499 : Address_next<= 61 ;
          500 : Address_next<= 30 ;
          502 : Address_next<= 31 ;
          503 : Address_next<= 62 ;
          504 : Address_next<= 124 ;
          506 : Address_next<= 125 ;
          507 : Address_next<= 62 ;
          509 : Address_next<= 63 ;
          510 : Address_next<= 126 ;
          512 : Address_next<= 127 ;
          513 : Address_next<= 63 ;
          514 : Address_next<= 31 ;
          515 : Address_next<= 15 ;
          516 : Address_next<= 7 ;
          517 : Address_next<= 3 ;
          518 : Address_next<= 1 ;
          525 : Address_next<= 1 ;
          526 : Address_next<= 1 ;
          527 : Address_next<= 2 ;
          528 : Address_next<= 4 ;
          529 : Address_next<= 8 ;
          530 : Address_next<= 16 ;
          531 : Address_next<= 32 ;
          532 : Address_next<= 64 ;
          533 : Address_next<= 128 ;
          535 : Address_next<= 129 ;
          536 : Address_next<= 64 ;
          538 : Address_next<= 65 ;
          539 : Address_next<= 130 ;
          541 : Address_next<= 131 ;
          542 : Address_next<= 65 ;
          543 : Address_next<= 32 ;
          545 : Address_next<= 33 ;
          546 : Address_next<= 66 ;
          547 : Address_next<= 132 ;
          549 : Address_next<= 133 ;
          550 : Address_next<= 66 ;
          552 : Address_next<= 67 ;
          553 : Address_next<= 134 ;
          555 : Address_next<= 135 ;
          556 : Address_next<= 67 ;
          557 : Address_next<= 33 ;
          558 : Address_next<= 16 ;
          560 : Address_next<= 17 ;
          561 : Address_next<= 34 ;
          562 : Address_next<= 68 ;
          563 : Address_next<= 136 ;
          565 : Address_next<= 137 ;
          566 : Address_next<= 68 ;
          568 : Address_next<= 69 ;
          569 : Address_next<= 138 ;
          571 : Address_next<= 139 ;
          572 : Address_next<= 69 ;
          573 : Address_next<= 34 ;
          575 : Address_next<= 35 ;
          576 : Address_next<= 70 ;
          577 : Address_next<= 140 ;
          579 : Address_next<= 141 ;
          580 : Address_next<= 70 ;
          582 : Address_next<= 71 ;
          583 : Address_next<= 142 ;
          585 : Address_next<= 143 ;
          586 : Address_next<= 71 ;
          587 : Address_next<= 35 ;
          588 : Address_next<= 17 ;
          589 : Address_next<= 8 ;
          591 : Address_next<= 9 ;
          592 : Address_next<= 18 ;
          593 : Address_next<= 36 ;
          594 : Address_next<= 72 ;
          595 : Address_next<= 144 ;
          597 : Address_next<= 145 ;
          598 : Address_next<= 72 ;
          600 : Address_next<= 73 ;
          601 : Address_next<= 146 ;
          603 : Address_next<= 147 ;
          604 : Address_next<= 73 ;
          605 : Address_next<= 36 ;
          607 : Address_next<= 37 ;
          608 : Address_next<= 74 ;
          609 : Address_next<= 148 ;
          611 : Address_next<= 149 ;
          612 : Address_next<= 74 ;
          614 : Address_next<= 75 ;
          615 : Address_next<= 150 ;
          617 : Address_next<= 151 ;
          618 : Address_next<= 75 ;
          619 : Address_next<= 37 ;
          620 : Address_next<= 18 ;
          622 : Address_next<= 19 ;
          623 : Address_next<= 38 ;
          624 : Address_next<= 76 ;
          625 : Address_next<= 152 ;
          627 : Address_next<= 153 ;
          628 : Address_next<= 76 ;
          630 : Address_next<= 77 ;
          631 : Address_next<= 154 ;
          633 : Address_next<= 155 ;
          634 : Address_next<= 77 ;
          635 : Address_next<= 38 ;
          637 : Address_next<= 39 ;
          638 : Address_next<= 78 ;
          639 : Address_next<= 156 ;
          641 : Address_next<= 157 ;
          642 : Address_next<= 78 ;
          644 : Address_next<= 79 ;
          645 : Address_next<= 158 ;
          647 : Address_next<= 159 ;
          648 : Address_next<= 79 ;
          649 : Address_next<= 39 ;
          650 : Address_next<= 19 ;
          651 : Address_next<= 9 ;
          652 : Address_next<= 4 ;
          654 : Address_next<= 5 ;
          655 : Address_next<= 10 ;
          656 : Address_next<= 20 ;
          657 : Address_next<= 40 ;
          658 : Address_next<= 80 ;
          659 : Address_next<= 160 ;
          661 : Address_next<= 161 ;
          662 : Address_next<= 80 ;
          664 : Address_next<= 81 ;
          665 : Address_next<= 162 ;
          667 : Address_next<= 163 ;
          668 : Address_next<= 81 ;
          669 : Address_next<= 40 ;
          671 : Address_next<= 41 ;
          672 : Address_next<= 82 ;
          673 : Address_next<= 164 ;
          675 : Address_next<= 165 ;
          676 : Address_next<= 82 ;
          678 : Address_next<= 83 ;
          679 : Address_next<= 166 ;
          681 : Address_next<= 167 ;
          682 : Address_next<= 83 ;
          683 : Address_next<= 41 ;
          684 : Address_next<= 20 ;
          686 : Address_next<= 21 ;
          687 : Address_next<= 42 ;
          688 : Address_next<= 84 ;
          689 : Address_next<= 168 ;
          691 : Address_next<= 169 ;
          692 : Address_next<= 84 ;
          694 : Address_next<= 85 ;
          695 : Address_next<= 170 ;
          697 : Address_next<= 171 ;
          698 : Address_next<= 85 ;
          699 : Address_next<= 42 ;
          701 : Address_next<= 43 ;
          702 : Address_next<= 86 ;
          703 : Address_next<= 172 ;
          705 : Address_next<= 173 ;
          706 : Address_next<= 86 ;
          708 : Address_next<= 87 ;
          709 : Address_next<= 174 ;
          711 : Address_next<= 175 ;
          712 : Address_next<= 87 ;
          713 : Address_next<= 43 ;
          714 : Address_next<= 21 ;
          715 : Address_next<= 10 ;
          717 : Address_next<= 11 ;
          718 : Address_next<= 22 ;
          719 : Address_next<= 44 ;
          720 : Address_next<= 88 ;
          721 : Address_next<= 176 ;
          723 : Address_next<= 177 ;
          724 : Address_next<= 88 ;
          726 : Address_next<= 89 ;
          727 : Address_next<= 178 ;
          729 : Address_next<= 179 ;
          730 : Address_next<= 89 ;
          731 : Address_next<= 44 ;
          733 : Address_next<= 45 ;
          734 : Address_next<= 90 ;
          735 : Address_next<= 180 ;
          737 : Address_next<= 181 ;
          738 : Address_next<= 90 ;
          740 : Address_next<= 91 ;
          741 : Address_next<= 182 ;
          743 : Address_next<= 183 ;
          744 : Address_next<= 91 ;
          745 : Address_next<= 45 ;
          746 : Address_next<= 22 ;
          748 : Address_next<= 23 ;
          749 : Address_next<= 46 ;
          750 : Address_next<= 92 ;
          751 : Address_next<= 184 ;
          753 : Address_next<= 185 ;
          754 : Address_next<= 92 ;
          756 : Address_next<= 93 ;
          757 : Address_next<= 186 ;
          759 : Address_next<= 187 ;
          760 : Address_next<= 93 ;
          761 : Address_next<= 46 ;
          763 : Address_next<= 47 ;
          764 : Address_next<= 94 ;
          765 : Address_next<= 188 ;
          767 : Address_next<= 189 ;
          768 : Address_next<= 94 ;
          770 : Address_next<= 95 ;
          771 : Address_next<= 190 ;
          773 : Address_next<= 191 ;
          774 : Address_next<= 95 ;
          775 : Address_next<= 47 ;
          776 : Address_next<= 23 ;
          777 : Address_next<= 11 ;
          778 : Address_next<= 5 ;
          779 : Address_next<= 2 ;
          782 : Address_next<= 3 ;
          783 : Address_next<= 6 ;
          784 : Address_next<= 12 ;
          785 : Address_next<= 24 ;
          786 : Address_next<= 48 ;
          787 : Address_next<= 96 ;
          788 : Address_next<= 192 ;
          790 : Address_next<= 193 ;
          791 : Address_next<= 96 ;
          793 : Address_next<= 97 ;
          794 : Address_next<= 194 ;
          796 : Address_next<= 195 ;
          797 : Address_next<= 97 ;
          798 : Address_next<= 48 ;
          800 : Address_next<= 49 ;
          801 : Address_next<= 98 ;
          802 : Address_next<= 196 ;
          804 : Address_next<= 197 ;
          805 : Address_next<= 98 ;
          807 : Address_next<= 99 ;
          808 : Address_next<= 198 ;
          810 : Address_next<= 199 ;
          811 : Address_next<= 99 ;
          812 : Address_next<= 49 ;
          813 : Address_next<= 24 ;
          815 : Address_next<= 25 ;
          816 : Address_next<= 50 ;
          817 : Address_next<= 100 ;
          818 : Address_next<= 200 ;
          820 : Address_next<= 201 ;
          821 : Address_next<= 100 ;
          823 : Address_next<= 101 ;
          824 : Address_next<= 202 ;
          826 : Address_next<= 203 ;
          827 : Address_next<= 101 ;
          828 : Address_next<= 50 ;
          830 : Address_next<= 51 ;
          831 : Address_next<= 102 ;
          832 : Address_next<= 204 ;
          834 : Address_next<= 205 ;
          835 : Address_next<= 102 ;
          837 : Address_next<= 103 ;
          838 : Address_next<= 206 ;
          840 : Address_next<= 207 ;
          841 : Address_next<= 103 ;
          842 : Address_next<= 51 ;
          843 : Address_next<= 25 ;
          844 : Address_next<= 12 ;
          846 : Address_next<= 13 ;
          847 : Address_next<= 26 ;
          848 : Address_next<= 52 ;
          849 : Address_next<= 104 ;
          850 : Address_next<= 208 ;
          852 : Address_next<= 209 ;
          853 : Address_next<= 104 ;
          855 : Address_next<= 105 ;
          856 : Address_next<= 210 ;
          858 : Address_next<= 211 ;
          859 : Address_next<= 105 ;
          860 : Address_next<= 52 ;
          862 : Address_next<= 53 ;
          863 : Address_next<= 106 ;
          864 : Address_next<= 212 ;
          866 : Address_next<= 213 ;
          867 : Address_next<= 106 ;
          869 : Address_next<= 107 ;
          870 : Address_next<= 214 ;
          872 : Address_next<= 215 ;
          873 : Address_next<= 107 ;
          874 : Address_next<= 53 ;
          875 : Address_next<= 26 ;
          877 : Address_next<= 27 ;
          878 : Address_next<= 54 ;
          879 : Address_next<= 108 ;
          880 : Address_next<= 216 ;
          882 : Address_next<= 217 ;
          883 : Address_next<= 108 ;
          885 : Address_next<= 109 ;
          886 : Address_next<= 218 ;
          888 : Address_next<= 219 ;
          889 : Address_next<= 109 ;
          890 : Address_next<= 54 ;
          892 : Address_next<= 55 ;
          893 : Address_next<= 110 ;
          894 : Address_next<= 220 ;
          896 : Address_next<= 221 ;
          897 : Address_next<= 110 ;
          899 : Address_next<= 111 ;
          900 : Address_next<= 222 ;
          902 : Address_next<= 223 ;
          903 : Address_next<= 111 ;
          904 : Address_next<= 55 ;
          905 : Address_next<= 27 ;
          906 : Address_next<= 13 ;
          907 : Address_next<= 6 ;
          909 : Address_next<= 7 ;
          910 : Address_next<= 14 ;
          911 : Address_next<= 28 ;
          912 : Address_next<= 56 ;
          913 : Address_next<= 112 ;
          914 : Address_next<= 224 ;
          916 : Address_next<= 225 ;
          917 : Address_next<= 112 ;
          919 : Address_next<= 113 ;
          920 : Address_next<= 226 ;
          922 : Address_next<= 227 ;
          923 : Address_next<= 113 ;
          924 : Address_next<= 56 ;
          926 : Address_next<= 57 ;
          927 : Address_next<= 114 ;
          928 : Address_next<= 228 ;
          930 : Address_next<= 229 ;
          931 : Address_next<= 114 ;
          933 : Address_next<= 115 ;
          934 : Address_next<= 230 ;
          936 : Address_next<= 231 ;
          937 : Address_next<= 115 ;
          938 : Address_next<= 57 ;
          939 : Address_next<= 28 ;
          941 : Address_next<= 29 ;
          942 : Address_next<= 58 ;
          943 : Address_next<= 116 ;
          944 : Address_next<= 232 ;
          946 : Address_next<= 233 ;
          947 : Address_next<= 116 ;
          949 : Address_next<= 117 ;
          950 : Address_next<= 234 ;
          952 : Address_next<= 235 ;
          953 : Address_next<= 117 ;
          954 : Address_next<= 58 ;
          956 : Address_next<= 59 ;
          957 : Address_next<= 118 ;
          958 : Address_next<= 236 ;
          960 : Address_next<= 237 ;
          961 : Address_next<= 118 ;
          963 : Address_next<= 119 ;
          964 : Address_next<= 238 ;
          966 : Address_next<= 239 ;
          967 : Address_next<= 119 ;
          968 : Address_next<= 59 ;
          969 : Address_next<= 29 ;
          970 : Address_next<= 14 ;
          972 : Address_next<= 15 ;
          973 : Address_next<= 30 ;
          974 : Address_next<= 60 ;
          975 : Address_next<= 120 ;
          976 : Address_next<= 240 ;
          978 : Address_next<= 241 ;
          979 : Address_next<= 120 ;
          981 : Address_next<= 121 ;
          982 : Address_next<= 242 ;
          984 : Address_next<= 243 ;
          985 : Address_next<= 121 ;
          986 : Address_next<= 60 ;
          988 : Address_next<= 61 ;
          989 : Address_next<= 122 ;
          990 : Address_next<= 244 ;
          992 : Address_next<= 245 ;
          993 : Address_next<= 122 ;
          995 : Address_next<= 123 ;
          996 : Address_next<= 246 ;
          998 : Address_next<= 247 ;
          999 : Address_next<= 123 ;
          1000 : Address_next<= 61 ;
          1001 : Address_next<= 30 ;
          1003 : Address_next<= 31 ;
          1004 : Address_next<= 62 ;
          1005 : Address_next<= 124 ;
          1006 : Address_next<= 248 ;
          1008 : Address_next<= 249 ;
          1009 : Address_next<= 124 ;
          1011 : Address_next<= 125 ;
          1012 : Address_next<= 250 ;
          1014 : Address_next<= 251 ;
          1015 : Address_next<= 125 ;
          1016 : Address_next<= 62 ;
          1018 : Address_next<= 63 ;
          1019 : Address_next<= 126 ;
          1020 : Address_next<= 252 ;
          1022 : Address_next<= 253 ;
          1023 : Address_next<= 126 ;
          1025 : Address_next<= 127 ;
          1026 : Address_next<= 254 ;
          1028 : Address_next<= 255 ;
          1029 : Address_next<= 127 ;
          1030 : Address_next<= 63 ;
          1031 : Address_next<= 31 ;
          1032 : Address_next<= 15 ;
          1033 : Address_next<= 7 ;
          1034 : Address_next<= 3 ;
          1035 : Address_next<= 1 ;
          1036 : Address_next<= 1 ;
          1049 : Address_next<= 1 ;
          1050 : Address_next<= 1 ;
          1051 : Address_next<= 1 ;
          1052 : Address_next<= 1 ;
          1053 : Address_next<= 2 ;
          1054 : Address_next<= 2 ;
          1055 : Address_next<= 4 ;
          1056 : Address_next<= 8 ;
          1057 : Address_next<= 16 ;
          1058 : Address_next<= 32 ;
          1059 : Address_next<= 64 ;
          1060 : Address_next<= 128 ;
          1061 : Address_next<= 256 ;
          1063 : Address_next<= 257 ;
          1064 : Address_next<= 128 ;
          1066 : Address_next<= 129 ;
          1067 : Address_next<= 258 ;
          1069 : Address_next<= 259 ;
          1070 : Address_next<= 129 ;
          1071 : Address_next<= 64 ;
          1073 : Address_next<= 65 ;
          1074 : Address_next<= 130 ;
          1075 : Address_next<= 260 ;
          1077 : Address_next<= 261 ;
          1078 : Address_next<= 130 ;
          1080 : Address_next<= 131 ;
          1081 : Address_next<= 262 ;
          1083 : Address_next<= 263 ;
          1084 : Address_next<= 131 ;
          1085 : Address_next<= 65 ;
          1086 : Address_next<= 32 ;
          1088 : Address_next<= 33 ;
          1089 : Address_next<= 66 ;
          1090 : Address_next<= 132 ;
          1091 : Address_next<= 264 ;
          1093 : Address_next<= 265 ;
          1094 : Address_next<= 132 ;
          1096 : Address_next<= 133 ;
          1097 : Address_next<= 266 ;
          1099 : Address_next<= 267 ;
          1100 : Address_next<= 133 ;
          1101 : Address_next<= 66 ;
          1103 : Address_next<= 67 ;
          1104 : Address_next<= 134 ;
          1105 : Address_next<= 268 ;
          1107 : Address_next<= 269 ;
          1108 : Address_next<= 134 ;
          1110 : Address_next<= 135 ;
          1111 : Address_next<= 270 ;
          1113 : Address_next<= 271 ;
          1114 : Address_next<= 135 ;
          1115 : Address_next<= 67 ;
          1116 : Address_next<= 33 ;
          1117 : Address_next<= 16 ;
          1119 : Address_next<= 17 ;
          1120 : Address_next<= 34 ;
          1121 : Address_next<= 68 ;
          1122 : Address_next<= 136 ;
          1123 : Address_next<= 272 ;
          1125 : Address_next<= 273 ;
          1126 : Address_next<= 136 ;
          1128 : Address_next<= 137 ;
          1129 : Address_next<= 274 ;
          1131 : Address_next<= 275 ;
          1132 : Address_next<= 137 ;
          1133 : Address_next<= 68 ;
          1135 : Address_next<= 69 ;
          1136 : Address_next<= 138 ;
          1137 : Address_next<= 276 ;
          1139 : Address_next<= 277 ;
          1140 : Address_next<= 138 ;
          1142 : Address_next<= 139 ;
          1143 : Address_next<= 278 ;
          1145 : Address_next<= 279 ;
          1146 : Address_next<= 139 ;
          1147 : Address_next<= 69 ;
          1148 : Address_next<= 34 ;
          1150 : Address_next<= 35 ;
          1151 : Address_next<= 70 ;
          1152 : Address_next<= 140 ;
          1153 : Address_next<= 280 ;
          1155 : Address_next<= 281 ;
          1156 : Address_next<= 140 ;
          1158 : Address_next<= 141 ;
          1159 : Address_next<= 282 ;
          1161 : Address_next<= 283 ;
          1162 : Address_next<= 141 ;
          1163 : Address_next<= 70 ;
          1165 : Address_next<= 71 ;
          1166 : Address_next<= 142 ;
          1167 : Address_next<= 284 ;
          1169 : Address_next<= 285 ;
          1170 : Address_next<= 142 ;
          1172 : Address_next<= 143 ;
          1173 : Address_next<= 286 ;
          1175 : Address_next<= 287 ;
          1176 : Address_next<= 143 ;
          1177 : Address_next<= 71 ;
          1178 : Address_next<= 35 ;
          1179 : Address_next<= 17 ;
          1180 : Address_next<= 8 ;
          1182 : Address_next<= 9 ;
          1183 : Address_next<= 18 ;
          1184 : Address_next<= 36 ;
          1185 : Address_next<= 72 ;
          1186 : Address_next<= 144 ;
          1187 : Address_next<= 288 ;
          1189 : Address_next<= 289 ;
          1190 : Address_next<= 144 ;
          1192 : Address_next<= 145 ;
          1193 : Address_next<= 290 ;
          1195 : Address_next<= 291 ;
          1196 : Address_next<= 145 ;
          1197 : Address_next<= 72 ;
          1199 : Address_next<= 73 ;
          1200 : Address_next<= 146 ;
          1201 : Address_next<= 292 ;
          1203 : Address_next<= 293 ;
          1204 : Address_next<= 146 ;
          1206 : Address_next<= 147 ;
          1207 : Address_next<= 294 ;
          1209 : Address_next<= 295 ;
          1210 : Address_next<= 147 ;
          1211 : Address_next<= 73 ;
          1212 : Address_next<= 36 ;
          1214 : Address_next<= 37 ;
          1215 : Address_next<= 74 ;
          1216 : Address_next<= 148 ;
          1217 : Address_next<= 296 ;
          1219 : Address_next<= 297 ;
          1220 : Address_next<= 148 ;
          1222 : Address_next<= 149 ;
          1223 : Address_next<= 298 ;
          1225 : Address_next<= 299 ;
          1226 : Address_next<= 149 ;
          1227 : Address_next<= 74 ;
          1229 : Address_next<= 75 ;
          1230 : Address_next<= 150 ;
          1231 : Address_next<= 300 ;
          1233 : Address_next<= 301 ;
          1234 : Address_next<= 150 ;
          1236 : Address_next<= 151 ;
          1237 : Address_next<= 302 ;
          1239 : Address_next<= 303 ;
          1240 : Address_next<= 151 ;
          1241 : Address_next<= 75 ;
          1242 : Address_next<= 37 ;
          1243 : Address_next<= 18 ;
          1245 : Address_next<= 19 ;
          1246 : Address_next<= 38 ;
          1247 : Address_next<= 76 ;
          1248 : Address_next<= 152 ;
          1249 : Address_next<= 304 ;
          1251 : Address_next<= 305 ;
          1252 : Address_next<= 152 ;
          1254 : Address_next<= 153 ;
          1255 : Address_next<= 306 ;
          1257 : Address_next<= 307 ;
          1258 : Address_next<= 153 ;
          1259 : Address_next<= 76 ;
          1261 : Address_next<= 77 ;
          1262 : Address_next<= 154 ;
          1263 : Address_next<= 308 ;
          1265 : Address_next<= 309 ;
          1266 : Address_next<= 154 ;
          1268 : Address_next<= 155 ;
          1269 : Address_next<= 310 ;
          1271 : Address_next<= 311 ;
          1272 : Address_next<= 155 ;
          1273 : Address_next<= 77 ;
          1274 : Address_next<= 38 ;
          1276 : Address_next<= 39 ;
          1277 : Address_next<= 78 ;
          1278 : Address_next<= 156 ;
          1279 : Address_next<= 312 ;
          1281 : Address_next<= 313 ;
          1282 : Address_next<= 156 ;
          1284 : Address_next<= 157 ;
          1285 : Address_next<= 314 ;
          1287 : Address_next<= 315 ;
          1288 : Address_next<= 157 ;
          1289 : Address_next<= 78 ;
          1291 : Address_next<= 79 ;
          1292 : Address_next<= 158 ;
          1293 : Address_next<= 316 ;
          1295 : Address_next<= 317 ;
          1296 : Address_next<= 158 ;
          1298 : Address_next<= 159 ;
          1299 : Address_next<= 318 ;
          1301 : Address_next<= 319 ;
          1302 : Address_next<= 159 ;
          1303 : Address_next<= 79 ;
          1304 : Address_next<= 39 ;
          1305 : Address_next<= 19 ;
          1306 : Address_next<= 9 ;
          1307 : Address_next<= 4 ;
          1310 : Address_next<= 5 ;
          1311 : Address_next<= 10 ;
          1312 : Address_next<= 20 ;
          1313 : Address_next<= 40 ;
          1314 : Address_next<= 80 ;
          1315 : Address_next<= 160 ;
          1316 : Address_next<= 320 ;
          1318 : Address_next<= 321 ;
          1319 : Address_next<= 160 ;
          1321 : Address_next<= 161 ;
          1322 : Address_next<= 322 ;
          1324 : Address_next<= 323 ;
          1325 : Address_next<= 161 ;
          1326 : Address_next<= 80 ;
          1328 : Address_next<= 81 ;
          1329 : Address_next<= 162 ;
          1330 : Address_next<= 324 ;
          1332 : Address_next<= 325 ;
          1333 : Address_next<= 162 ;
          1335 : Address_next<= 163 ;
          1336 : Address_next<= 326 ;
          1338 : Address_next<= 327 ;
          1339 : Address_next<= 163 ;
          1340 : Address_next<= 81 ;
          1341 : Address_next<= 40 ;
          1343 : Address_next<= 41 ;
          1344 : Address_next<= 82 ;
          1345 : Address_next<= 164 ;
          1346 : Address_next<= 328 ;
          1348 : Address_next<= 329 ;
          1349 : Address_next<= 164 ;
          1351 : Address_next<= 165 ;
          1352 : Address_next<= 330 ;
          1354 : Address_next<= 331 ;
          1355 : Address_next<= 165 ;
          1356 : Address_next<= 82 ;
          1358 : Address_next<= 83 ;
          1359 : Address_next<= 166 ;
          1360 : Address_next<= 332 ;
          1362 : Address_next<= 333 ;
          1363 : Address_next<= 166 ;
          1365 : Address_next<= 167 ;
          1366 : Address_next<= 334 ;
          1368 : Address_next<= 335 ;
          1369 : Address_next<= 167 ;
          1370 : Address_next<= 83 ;
          1371 : Address_next<= 41 ;
          1372 : Address_next<= 20 ;
          1374 : Address_next<= 21 ;
          1375 : Address_next<= 42 ;
          1376 : Address_next<= 84 ;
          1377 : Address_next<= 168 ;
          1378 : Address_next<= 336 ;
          1380 : Address_next<= 337 ;
          1381 : Address_next<= 168 ;
          1383 : Address_next<= 169 ;
          1384 : Address_next<= 338 ;
          1386 : Address_next<= 339 ;
          1387 : Address_next<= 169 ;
          1388 : Address_next<= 84 ;
          1390 : Address_next<= 85 ;
          1391 : Address_next<= 170 ;
          1392 : Address_next<= 340 ;
          1394 : Address_next<= 341 ;
          1395 : Address_next<= 170 ;
          1397 : Address_next<= 171 ;
          1398 : Address_next<= 342 ;
          1400 : Address_next<= 343 ;
          1401 : Address_next<= 171 ;
          1402 : Address_next<= 85 ;
          1403 : Address_next<= 42 ;
          1405 : Address_next<= 43 ;
          1406 : Address_next<= 86 ;
          1407 : Address_next<= 172 ;
          1408 : Address_next<= 344 ;
          1410 : Address_next<= 345 ;
          1411 : Address_next<= 172 ;
          1413 : Address_next<= 173 ;
          1414 : Address_next<= 346 ;
          1416 : Address_next<= 347 ;
          1417 : Address_next<= 173 ;
          1418 : Address_next<= 86 ;
          1420 : Address_next<= 87 ;
          1421 : Address_next<= 174 ;
          1422 : Address_next<= 348 ;
          1424 : Address_next<= 349 ;
          1425 : Address_next<= 174 ;
          1427 : Address_next<= 175 ;
          1428 : Address_next<= 350 ;
          1430 : Address_next<= 351 ;
          1431 : Address_next<= 175 ;
          1432 : Address_next<= 87 ;
          1433 : Address_next<= 43 ;
          1434 : Address_next<= 21 ;
          1435 : Address_next<= 10 ;
          1437 : Address_next<= 11 ;
          1438 : Address_next<= 22 ;
          1439 : Address_next<= 44 ;
          1440 : Address_next<= 88 ;
          1441 : Address_next<= 176 ;
          1442 : Address_next<= 352 ;
          1444 : Address_next<= 353 ;
          1445 : Address_next<= 176 ;
          1447 : Address_next<= 177 ;
          1448 : Address_next<= 354 ;
          1450 : Address_next<= 355 ;
          1451 : Address_next<= 177 ;
          1452 : Address_next<= 88 ;
          1454 : Address_next<= 89 ;
          1455 : Address_next<= 178 ;
          1456 : Address_next<= 356 ;
          1458 : Address_next<= 357 ;
          1459 : Address_next<= 178 ;
          1461 : Address_next<= 179 ;
          1462 : Address_next<= 358 ;
          1464 : Address_next<= 359 ;
          1465 : Address_next<= 179 ;
          1466 : Address_next<= 89 ;
          1467 : Address_next<= 44 ;
          1469 : Address_next<= 45 ;
          1470 : Address_next<= 90 ;
          1471 : Address_next<= 180 ;
          1472 : Address_next<= 360 ;
          1474 : Address_next<= 361 ;
          1475 : Address_next<= 180 ;
          1477 : Address_next<= 181 ;
          1478 : Address_next<= 362 ;
          1480 : Address_next<= 363 ;
          1481 : Address_next<= 181 ;
          1482 : Address_next<= 90 ;
          1484 : Address_next<= 91 ;
          1485 : Address_next<= 182 ;
          1486 : Address_next<= 364 ;
          1488 : Address_next<= 365 ;
          1489 : Address_next<= 182 ;
          1491 : Address_next<= 183 ;
          1492 : Address_next<= 366 ;
          1494 : Address_next<= 367 ;
          1495 : Address_next<= 183 ;
          1496 : Address_next<= 91 ;
          1497 : Address_next<= 45 ;
          1498 : Address_next<= 22 ;
          1500 : Address_next<= 23 ;
          1501 : Address_next<= 46 ;
          1502 : Address_next<= 92 ;
          1503 : Address_next<= 184 ;
          1504 : Address_next<= 368 ;
          1506 : Address_next<= 369 ;
          1507 : Address_next<= 184 ;
          1509 : Address_next<= 185 ;
          1510 : Address_next<= 370 ;
          1512 : Address_next<= 371 ;
          1513 : Address_next<= 185 ;
          1514 : Address_next<= 92 ;
          1516 : Address_next<= 93 ;
          1517 : Address_next<= 186 ;
          1518 : Address_next<= 372 ;
          1520 : Address_next<= 373 ;
          1521 : Address_next<= 186 ;
          1523 : Address_next<= 187 ;
          1524 : Address_next<= 374 ;
          1526 : Address_next<= 375 ;
          1527 : Address_next<= 187 ;
          1528 : Address_next<= 93 ;
          1529 : Address_next<= 46 ;
          1531 : Address_next<= 47 ;
          1532 : Address_next<= 94 ;
          1533 : Address_next<= 188 ;
          1534 : Address_next<= 376 ;
          1536 : Address_next<= 377 ;
          1537 : Address_next<= 188 ;
          1539 : Address_next<= 189 ;
          1540 : Address_next<= 378 ;
          1542 : Address_next<= 379 ;
          1543 : Address_next<= 189 ;
          1544 : Address_next<= 94 ;
          1546 : Address_next<= 95 ;
          1547 : Address_next<= 190 ;
          1548 : Address_next<= 380 ;
          1550 : Address_next<= 381 ;
          1551 : Address_next<= 190 ;
          1553 : Address_next<= 191 ;
          1554 : Address_next<= 382 ;
          1556 : Address_next<= 383 ;
          1557 : Address_next<= 191 ;
          1558 : Address_next<= 95 ;
          1559 : Address_next<= 47 ;
          1560 : Address_next<= 23 ;
          1561 : Address_next<= 11 ;
          1562 : Address_next<= 5 ;
          1563 : Address_next<= 2 ;
          1564 : Address_next<= 2 ;
          1569 : Address_next<= 3 ;
          1570 : Address_next<= 3 ;
          1571 : Address_next<= 6 ;
          1572 : Address_next<= 12 ;
          1573 : Address_next<= 24 ;
          1574 : Address_next<= 48 ;
          1575 : Address_next<= 96 ;
          1576 : Address_next<= 192 ;
          1577 : Address_next<= 384 ;
          1579 : Address_next<= 385 ;
          1580 : Address_next<= 192 ;
          1582 : Address_next<= 193 ;
          1583 : Address_next<= 386 ;
          1585 : Address_next<= 387 ;
          1586 : Address_next<= 193 ;
          1587 : Address_next<= 96 ;
          1589 : Address_next<= 97 ;
          1590 : Address_next<= 194 ;
          1591 : Address_next<= 388 ;
          1593 : Address_next<= 389 ;
          1594 : Address_next<= 194 ;
          1596 : Address_next<= 195 ;
          1597 : Address_next<= 390 ;
          1599 : Address_next<= 391 ;
          1600 : Address_next<= 195 ;
          1601 : Address_next<= 97 ;
          1602 : Address_next<= 48 ;
          1604 : Address_next<= 49 ;
          1605 : Address_next<= 98 ;
          1606 : Address_next<= 196 ;
          1607 : Address_next<= 392 ;
          1609 : Address_next<= 393 ;
          1610 : Address_next<= 196 ;
          1612 : Address_next<= 197 ;
          1613 : Address_next<= 394 ;
          1615 : Address_next<= 395 ;
          1616 : Address_next<= 197 ;
          1617 : Address_next<= 98 ;
          1619 : Address_next<= 99 ;
          1620 : Address_next<= 198 ;
          1621 : Address_next<= 396 ;
          1623 : Address_next<= 397 ;
          1624 : Address_next<= 198 ;
          1626 : Address_next<= 199 ;
          1627 : Address_next<= 398 ;
          1629 : Address_next<= 399 ;
          1630 : Address_next<= 199 ;
          1631 : Address_next<= 99 ;
          1632 : Address_next<= 49 ;
          1633 : Address_next<= 24 ;
          1635 : Address_next<= 25 ;
          1636 : Address_next<= 50 ;
          1637 : Address_next<= 100 ;
          1638 : Address_next<= 200 ;
          1639 : Address_next<= 400 ;
          1641 : Address_next<= 401 ;
          1642 : Address_next<= 200 ;
          1644 : Address_next<= 201 ;
          1645 : Address_next<= 402 ;
          1647 : Address_next<= 403 ;
          1648 : Address_next<= 201 ;
          1649 : Address_next<= 100 ;
          1651 : Address_next<= 101 ;
          1652 : Address_next<= 202 ;
          1653 : Address_next<= 404 ;
          1655 : Address_next<= 405 ;
          1656 : Address_next<= 202 ;
          1658 : Address_next<= 203 ;
          1659 : Address_next<= 406 ;
          1661 : Address_next<= 407 ;
          1662 : Address_next<= 203 ;
          1663 : Address_next<= 101 ;
          1664 : Address_next<= 50 ;
          1666 : Address_next<= 51 ;
          1667 : Address_next<= 102 ;
          1668 : Address_next<= 204 ;
          1669 : Address_next<= 408 ;
          1671 : Address_next<= 409 ;
          1672 : Address_next<= 204 ;
          1674 : Address_next<= 205 ;
          1675 : Address_next<= 410 ;
          1677 : Address_next<= 411 ;
          1678 : Address_next<= 205 ;
          1679 : Address_next<= 102 ;
          1681 : Address_next<= 103 ;
          1682 : Address_next<= 206 ;
          1683 : Address_next<= 412 ;
          1685 : Address_next<= 413 ;
          1686 : Address_next<= 206 ;
          1688 : Address_next<= 207 ;
          1689 : Address_next<= 414 ;
          1691 : Address_next<= 415 ;
          1692 : Address_next<= 207 ;
          1693 : Address_next<= 103 ;
          1694 : Address_next<= 51 ;
          1695 : Address_next<= 25 ;
          1696 : Address_next<= 12 ;
          1698 : Address_next<= 13 ;
          1699 : Address_next<= 26 ;
          1700 : Address_next<= 52 ;
          1701 : Address_next<= 104 ;
          1702 : Address_next<= 208 ;
          1703 : Address_next<= 416 ;
          1705 : Address_next<= 417 ;
          1706 : Address_next<= 208 ;
          1708 : Address_next<= 209 ;
          1709 : Address_next<= 418 ;
          1711 : Address_next<= 419 ;
          1712 : Address_next<= 209 ;
          1713 : Address_next<= 104 ;
          1715 : Address_next<= 105 ;
          1716 : Address_next<= 210 ;
          1717 : Address_next<= 420 ;
          1719 : Address_next<= 421 ;
          1720 : Address_next<= 210 ;
          1722 : Address_next<= 211 ;
          1723 : Address_next<= 422 ;
          1725 : Address_next<= 423 ;
          1726 : Address_next<= 211 ;
          1727 : Address_next<= 105 ;
          1728 : Address_next<= 52 ;
          1730 : Address_next<= 53 ;
          1731 : Address_next<= 106 ;
          1732 : Address_next<= 212 ;
          1733 : Address_next<= 424 ;
          1735 : Address_next<= 425 ;
          1736 : Address_next<= 212 ;
          1738 : Address_next<= 213 ;
          1739 : Address_next<= 426 ;
          1741 : Address_next<= 427 ;
          1742 : Address_next<= 213 ;
          1743 : Address_next<= 106 ;
          1745 : Address_next<= 107 ;
          1746 : Address_next<= 214 ;
          1747 : Address_next<= 428 ;
          1749 : Address_next<= 429 ;
          1750 : Address_next<= 214 ;
          1752 : Address_next<= 215 ;
          1753 : Address_next<= 430 ;
          1755 : Address_next<= 431 ;
          1756 : Address_next<= 215 ;
          1757 : Address_next<= 107 ;
          1758 : Address_next<= 53 ;
          1759 : Address_next<= 26 ;
          1761 : Address_next<= 27 ;
          1762 : Address_next<= 54 ;
          1763 : Address_next<= 108 ;
          1764 : Address_next<= 216 ;
          1765 : Address_next<= 432 ;
          1767 : Address_next<= 433 ;
          1768 : Address_next<= 216 ;
          1770 : Address_next<= 217 ;
          1771 : Address_next<= 434 ;
          1773 : Address_next<= 435 ;
          1774 : Address_next<= 217 ;
          1775 : Address_next<= 108 ;
          1777 : Address_next<= 109 ;
          1778 : Address_next<= 218 ;
          1779 : Address_next<= 436 ;
          1781 : Address_next<= 437 ;
          1782 : Address_next<= 218 ;
          1784 : Address_next<= 219 ;
          1785 : Address_next<= 438 ;
          1787 : Address_next<= 439 ;
          1788 : Address_next<= 219 ;
          1789 : Address_next<= 109 ;
          1790 : Address_next<= 54 ;
          1792 : Address_next<= 55 ;
          1793 : Address_next<= 110 ;
          1794 : Address_next<= 220 ;
          1795 : Address_next<= 440 ;
          1797 : Address_next<= 441 ;
          1798 : Address_next<= 220 ;
          1800 : Address_next<= 221 ;
          1801 : Address_next<= 442 ;
          1803 : Address_next<= 443 ;
          1804 : Address_next<= 221 ;
          1805 : Address_next<= 110 ;
          1807 : Address_next<= 111 ;
          1808 : Address_next<= 222 ;
          1809 : Address_next<= 444 ;
          1811 : Address_next<= 445 ;
          1812 : Address_next<= 222 ;
          1814 : Address_next<= 223 ;
          1815 : Address_next<= 446 ;
          1817 : Address_next<= 447 ;
          1818 : Address_next<= 223 ;
          1819 : Address_next<= 111 ;
          1820 : Address_next<= 55 ;
          1821 : Address_next<= 27 ;
          1822 : Address_next<= 13 ;
          1823 : Address_next<= 6 ;
          1826 : Address_next<= 7 ;
          1827 : Address_next<= 14 ;
          1828 : Address_next<= 28 ;
          1829 : Address_next<= 56 ;
          1830 : Address_next<= 112 ;
          1831 : Address_next<= 224 ;
          1832 : Address_next<= 448 ;
          1834 : Address_next<= 449 ;
          1835 : Address_next<= 224 ;
          1837 : Address_next<= 225 ;
          1838 : Address_next<= 450 ;
          1840 : Address_next<= 451 ;
          1841 : Address_next<= 225 ;
          1842 : Address_next<= 112 ;
          1844 : Address_next<= 113 ;
          1845 : Address_next<= 226 ;
          1846 : Address_next<= 452 ;
          1848 : Address_next<= 453 ;
          1849 : Address_next<= 226 ;
          1851 : Address_next<= 227 ;
          1852 : Address_next<= 454 ;
          1854 : Address_next<= 455 ;
          1855 : Address_next<= 227 ;
          1856 : Address_next<= 113 ;
          1857 : Address_next<= 56 ;
          1859 : Address_next<= 57 ;
          1860 : Address_next<= 114 ;
          1861 : Address_next<= 228 ;
          1862 : Address_next<= 456 ;
          1864 : Address_next<= 457 ;
          1865 : Address_next<= 228 ;
          1867 : Address_next<= 229 ;
          1868 : Address_next<= 458 ;
          1870 : Address_next<= 459 ;
          1871 : Address_next<= 229 ;
          1872 : Address_next<= 114 ;
          1874 : Address_next<= 115 ;
          1875 : Address_next<= 230 ;
          1876 : Address_next<= 460 ;
          1878 : Address_next<= 461 ;
          1879 : Address_next<= 230 ;
          1881 : Address_next<= 231 ;
          1882 : Address_next<= 462 ;
          1884 : Address_next<= 463 ;
          1885 : Address_next<= 231 ;
          1886 : Address_next<= 115 ;
          1887 : Address_next<= 57 ;
          1888 : Address_next<= 28 ;
          1890 : Address_next<= 29 ;
          1891 : Address_next<= 58 ;
          1892 : Address_next<= 116 ;
          1893 : Address_next<= 232 ;
          1894 : Address_next<= 464 ;
          1896 : Address_next<= 465 ;
          1897 : Address_next<= 232 ;
          1899 : Address_next<= 233 ;
          1900 : Address_next<= 466 ;
          1902 : Address_next<= 467 ;
          1903 : Address_next<= 233 ;
          1904 : Address_next<= 116 ;
          1906 : Address_next<= 117 ;
          1907 : Address_next<= 234 ;
          1908 : Address_next<= 468 ;
          1910 : Address_next<= 469 ;
          1911 : Address_next<= 234 ;
          1913 : Address_next<= 235 ;
          1914 : Address_next<= 470 ;
          1916 : Address_next<= 471 ;
          1917 : Address_next<= 235 ;
          1918 : Address_next<= 117 ;
          1919 : Address_next<= 58 ;
          1921 : Address_next<= 59 ;
          1922 : Address_next<= 118 ;
          1923 : Address_next<= 236 ;
          1924 : Address_next<= 472 ;
          1926 : Address_next<= 473 ;
          1927 : Address_next<= 236 ;
          1929 : Address_next<= 237 ;
          1930 : Address_next<= 474 ;
          1932 : Address_next<= 475 ;
          1933 : Address_next<= 237 ;
          1934 : Address_next<= 118 ;
          1936 : Address_next<= 119 ;
          1937 : Address_next<= 238 ;
          1938 : Address_next<= 476 ;
          1940 : Address_next<= 477 ;
          1941 : Address_next<= 238 ;
          1943 : Address_next<= 239 ;
          1944 : Address_next<= 478 ;
          1946 : Address_next<= 479 ;
          1947 : Address_next<= 239 ;
          1948 : Address_next<= 119 ;
          1949 : Address_next<= 59 ;
          1950 : Address_next<= 29 ;
          1951 : Address_next<= 14 ;
          1953 : Address_next<= 15 ;
          1954 : Address_next<= 30 ;
          1955 : Address_next<= 60 ;
          1956 : Address_next<= 120 ;
          1957 : Address_next<= 240 ;
          1958 : Address_next<= 480 ;
          1960 : Address_next<= 481 ;
          1961 : Address_next<= 240 ;
          1963 : Address_next<= 241 ;
          1964 : Address_next<= 482 ;
          1966 : Address_next<= 483 ;
          1967 : Address_next<= 241 ;
          1968 : Address_next<= 120 ;
          1970 : Address_next<= 121 ;
          1971 : Address_next<= 242 ;
          1972 : Address_next<= 484 ;
          1974 : Address_next<= 485 ;
          1975 : Address_next<= 242 ;
          1977 : Address_next<= 243 ;
          1978 : Address_next<= 486 ;
          1980 : Address_next<= 487 ;
          1981 : Address_next<= 243 ;
          1982 : Address_next<= 121 ;
          1983 : Address_next<= 60 ;
          1985 : Address_next<= 61 ;
          1986 : Address_next<= 122 ;
          1987 : Address_next<= 244 ;
          1988 : Address_next<= 488 ;
          1990 : Address_next<= 489 ;
          1991 : Address_next<= 244 ;
          1993 : Address_next<= 245 ;
          1994 : Address_next<= 490 ;
          1996 : Address_next<= 491 ;
          1997 : Address_next<= 245 ;
          1998 : Address_next<= 122 ;
          2000 : Address_next<= 123 ;
          2001 : Address_next<= 246 ;
          2002 : Address_next<= 492 ;
          2004 : Address_next<= 493 ;
          2005 : Address_next<= 246 ;
          2007 : Address_next<= 247 ;
          2008 : Address_next<= 494 ;
          2010 : Address_next<= 495 ;
          2011 : Address_next<= 247 ;
          2012 : Address_next<= 123 ;
          2013 : Address_next<= 61 ;
          2014 : Address_next<= 30 ;
          2016 : Address_next<= 31 ;
          2017 : Address_next<= 62 ;
          2018 : Address_next<= 124 ;
          2019 : Address_next<= 248 ;
          2020 : Address_next<= 496 ;
          2022 : Address_next<= 497 ;
          2023 : Address_next<= 248 ;
          2025 : Address_next<= 249 ;
          2026 : Address_next<= 498 ;
          2028 : Address_next<= 499 ;
          2029 : Address_next<= 249 ;
          2030 : Address_next<= 124 ;
          2032 : Address_next<= 125 ;
          2033 : Address_next<= 250 ;
          2034 : Address_next<= 500 ;
          2036 : Address_next<= 501 ;
          2037 : Address_next<= 250 ;
          2039 : Address_next<= 251 ;
          2040 : Address_next<= 502 ;
          2042 : Address_next<= 503 ;
          2043 : Address_next<= 251 ;
          2044 : Address_next<= 125 ;
          2045 : Address_next<= 62 ;
          2047 : Address_next<= 63 ;
          2048 : Address_next<= 126 ;
          2049 : Address_next<= 252 ;
          2050 : Address_next<= 504 ;
          2052 : Address_next<= 505 ;
          2053 : Address_next<= 252 ;
          2055 : Address_next<= 253 ;
          2056 : Address_next<= 506 ;
          2058 : Address_next<= 507 ;
          2059 : Address_next<= 253 ;
          2060 : Address_next<= 126 ;
          2062 : Address_next<= 127 ;
          2063 : Address_next<= 254 ;
          2064 : Address_next<= 508 ;
          2066 : Address_next<= 509 ;
          2067 : Address_next<= 254 ;
          2069 : Address_next<= 255 ;
          2070 : Address_next<= 510 ;
          2072 : Address_next<= 511 ;
          2073 : Address_next<= 255 ;
          2074 : Address_next<= 127 ;
          2075 : Address_next<= 63 ;
          2076 : Address_next<= 31 ;
          2077 : Address_next<= 15 ;
          2078 : Address_next<= 7 ;
          2079 : Address_next<= 3 ;
          2080 : Address_next<= 3 ;
          2081 : Address_next<= 1 ;
          2082 : Address_next<= 1 ;
          2083 : Address_next<= 1 ;
          2084 : Address_next<= 1 ;
       endcase


      end
      else begin
           L_Nv_next                     <=1024;
           L_opcode_next <= TYPE1;
           L_part_count_next <= 0;
           Address_next <= 0;
      end
end
end
endmodule


