module opcode #(parameter P = 16) (clk, rst, channel, I_program_counter,O_opcode, O_opcode_next, O_opcode_delay,
        O_Nv,O_Nv_next, O_part_count,O_part_count_next, O_address, O_address_next, O_opcode_before, O_Nv_before, O_bit_count);
        input clk,rst;
        input channel;
        input [15:0] I_program_counter;
        output [3:0] O_opcode,O_opcode_next, O_opcode_before, O_opcode_delay;
        output [10:0] O_Nv, O_Nv_next, O_Nv_before;
        output [5:0] O_part_count, O_part_count_next;
        output [9:0] O_address, O_address_next;
        output [12:0] O_bit_count;
        localparam TYPE1     = 4'b0000;
        localparam TYPE2     = 4'b0001;
        localparam BOTTOM    = 4'b0010;
        localparam TYPE3     = 4'b0011;
        localparam IDLE      = 4'b1011;

        reg [3:0] L_opcode, L_opcode_next, L_opcode_before, L_opcode_delay;
        reg [10:0] L_Nv,L_Nv_next,L_Nv_before, L_Nv_delay;
        reg [5:0] L_part_count, L_part_count_next, L_part_count_delay;
        reg [9:0] Address, Address_next, Address_delay;
        reg[12:0] L_bit_count;
        
        // assignment of outputs
        assign O_opcode = L_opcode;
        assign O_opcode_delay = L_opcode_delay;
        assign O_opcode_next = L_opcode_next;
        assign O_opcode_before = L_opcode_before;
        assign O_Nv = L_Nv;
        assign O_Nv_next = L_Nv_next;
        assign O_Nv_before = L_Nv_before;
        assign O_part_count = L_part_count;
        assign O_part_count_next = L_part_count_next;
        assign O_address = Address;
        assign O_address_next = Address_next;
        assign O_bit_count = L_bit_count;


        wire islast, oprand;
       assign islast = (L_Nv_next) > (2*P*(1+L_part_count_next));
       assign oprand = (L_opcode_next==TYPE1||L_opcode_next==TYPE2);

       always @(posedge clk)
     begin       
           if(!rst) begin
                L_Nv_before <= L_Nv;        
                L_Nv <= L_Nv_delay;
                L_Nv_delay <= L_Nv_next;

                L_opcode_before <= L_opcode;
                L_opcode <= L_opcode_delay;
                L_opcode_delay <= L_opcode_next;


                L_part_count <= L_part_count_delay;
                L_part_count_delay <= L_part_count_next;

//                Address_before <= Address;       
                L_bit_count <= (L_bit_count+2*(L_opcode==BOTTOM));

                Address <= Address_delay;
                Address_delay <= Address_next;
            end
            else begin
              L_bit_count <= 0;
              L_Nv                          <=1024; 
              L_Nv_before                          <=1024; 
              L_Nv_delay                          <=1024; 

              L_opcode_before <= TYPE1;
              L_opcode <= TYPE1;
              L_opcode_delay <= TYPE1;


              L_part_count <= 0;
              L_part_count_delay <= 0;

              Address <= 0;
              Address_delay <= 0;
            end
        end



        always @(posedge clk) begin
            if(rst) begin
            
            L_Nv_next                     <=1024;
            L_opcode_next <= TYPE1;
            L_part_count_next <= 0;
            // Address <= -1;
            Address_next <= 0;
            end
            else begin
           if (channel) begin
              case (L_Nv_next)
                1024 : L_Nv_next <= islast ? 1024 : 512;
                512 : L_Nv_next <= islast ?  512 : (oprand?256:1024);
                256 : L_Nv_next <= islast ? 256 : (oprand?128:512);
                128 : L_Nv_next <= oprand ? 64 : 256;
                64 : L_Nv_next <= oprand ? 32 : 128;
                32 : L_Nv_next <= oprand ? 16 : 64;
                16 : L_Nv_next <= oprand ? 8 : 32;
                8 : L_Nv_next <= oprand ? 4 : 16;
                4 : L_Nv_next <= oprand ? 2 : 8;
                2 : L_Nv_next <= 4;
                default: L_Nv_next <= 1024;
              endcase

              case (L_opcode_next)
                TYPE1 : L_opcode_next <= islast ? TYPE1 : ( (L_Nv_next==4) ? BOTTOM : TYPE1 );
                TYPE2 : L_opcode_next <= islast ? TYPE2 : ( (L_Nv_next==4) ? BOTTOM : TYPE1 );
                TYPE3 : L_opcode_next <= islast ? TYPE3 : ( (Address_next[0]) ? TYPE3 : TYPE2);
                BOTTOM : L_opcode_next <= Address_next[0] ? TYPE3 : TYPE2 ;
                default: L_opcode_next <= TYPE1;
              endcase

                // case (L_part_count_next)
                //   0 : L_part_count_next <= (L_Nv_next>2*P) ? 1 : 0;
                //   1 : L_part_count_next <= (L_Nv_next>4*P) ? 2 : 0;
                //   2 : L_part_count_next <= (L_Nv_next>4*P) ? 3 : 0;
                //   3 : L_part_count_next <=  0;
                //   4 : L_part_count_next <= (L_Nv_next>8*P) ? 5 : 0;
                //   5 : L_part_count_next <= (L_Nv_next>8*P) ? 6 : 0;
                //   6 : L_part_count_next <= (L_Nv_next>8*P) ? 7 : 0;
                //   7 : L_part_count_next <= 0;
                //   default: L_part_count_next <= 0;
                // endcase
                L_part_count_next <= islast ? (L_part_count_next+1) : 0;


          

       case(I_program_counter)
        65 : Address_next<= 1 ;
        68 : Address_next<= 1 ;
        69 : Address_next<= 2 ;
        71 : Address_next<= 3 ;
        72 : Address_next<= 1 ;
        75 : Address_next<= 1 ;
        76 : Address_next<= 2 ;
        77 : Address_next<= 4 ;
        79 : Address_next<= 5 ;
        80 : Address_next<= 2 ;
        82 : Address_next<= 3 ;
        83 : Address_next<= 6 ;
        85 : Address_next<= 7 ;
        86 : Address_next<= 3 ;
        87 : Address_next<= 1 ;
        90 : Address_next<= 1 ;
        91 : Address_next<= 2 ;
        92 : Address_next<= 4 ;
        93 : Address_next<= 8 ;
        95 : Address_next<= 9 ;
        96 : Address_next<= 4 ;
        98 : Address_next<= 5 ;
        99 : Address_next<= 10 ;
        101 : Address_next<= 11 ;
        102 : Address_next<= 5 ;
        103 : Address_next<= 2 ;
        105 : Address_next<= 3 ;
        106 : Address_next<= 6 ;
        107 : Address_next<= 12 ;
        109 : Address_next<= 13 ;
        110 : Address_next<= 6 ;
        112 : Address_next<= 7 ;
        113 : Address_next<= 14 ;
        115 : Address_next<= 15 ;
        116 : Address_next<= 7 ;
        117 : Address_next<= 3 ;
        118 : Address_next<= 1 ;
        122 : Address_next<= 1 ;
        123 : Address_next<= 2 ;
        124 : Address_next<= 4 ;
        125 : Address_next<= 8 ;
        126 : Address_next<= 16 ;
        128 : Address_next<= 17 ;
        129 : Address_next<= 8 ;
        131 : Address_next<= 9 ;
        132 : Address_next<= 18 ;
        134 : Address_next<= 19 ;
        135 : Address_next<= 9 ;
        136 : Address_next<= 4 ;
        138 : Address_next<= 5 ;
        139 : Address_next<= 10 ;
        140 : Address_next<= 20 ;
        142 : Address_next<= 21 ;
        143 : Address_next<= 10 ;
        145 : Address_next<= 11 ;
        146 : Address_next<= 22 ;
        148 : Address_next<= 23 ;
        149 : Address_next<= 11 ;
        150 : Address_next<= 5 ;
        151 : Address_next<= 2 ;
        153 : Address_next<= 3 ;
        154 : Address_next<= 6 ;
        155 : Address_next<= 12 ;
        156 : Address_next<= 24 ;
        158 : Address_next<= 25 ;
        159 : Address_next<= 12 ;
        161 : Address_next<= 13 ;
        162 : Address_next<= 26 ;
        164 : Address_next<= 27 ;
        165 : Address_next<= 13 ;
        166 : Address_next<= 6 ;
        168 : Address_next<= 7 ;
        169 : Address_next<= 14 ;
        170 : Address_next<= 28 ;
        172 : Address_next<= 29 ;
        173 : Address_next<= 14 ;
        175 : Address_next<= 15 ;
        176 : Address_next<= 30 ;
        178 : Address_next<= 31 ;
        179 : Address_next<= 15 ;
        180 : Address_next<= 7 ;
        181 : Address_next<= 3 ;
        182 : Address_next<= 1 ;
        189 : Address_next<= 1 ;
        190 : Address_next<= 1 ;
        191 : Address_next<= 2 ;
        192 : Address_next<= 4 ;
        193 : Address_next<= 8 ;
        194 : Address_next<= 16 ;
        195 : Address_next<= 32 ;
        197 : Address_next<= 33 ;
        198 : Address_next<= 16 ;
        200 : Address_next<= 17 ;
        201 : Address_next<= 34 ;
        203 : Address_next<= 35 ;
        204 : Address_next<= 17 ;
        205 : Address_next<= 8 ;
        207 : Address_next<= 9 ;
        208 : Address_next<= 18 ;
        209 : Address_next<= 36 ;
        211 : Address_next<= 37 ;
        212 : Address_next<= 18 ;
        214 : Address_next<= 19 ;
        215 : Address_next<= 38 ;
        217 : Address_next<= 39 ;
        218 : Address_next<= 19 ;
        219 : Address_next<= 9 ;
        220 : Address_next<= 4 ;
        222 : Address_next<= 5 ;
        223 : Address_next<= 10 ;
        224 : Address_next<= 20 ;
        225 : Address_next<= 40 ;
        227 : Address_next<= 41 ;
        228 : Address_next<= 20 ;
        230 : Address_next<= 21 ;
        231 : Address_next<= 42 ;
        233 : Address_next<= 43 ;
        234 : Address_next<= 21 ;
        235 : Address_next<= 10 ;
        237 : Address_next<= 11 ;
        238 : Address_next<= 22 ;
        239 : Address_next<= 44 ;
        241 : Address_next<= 45 ;
        242 : Address_next<= 22 ;
        244 : Address_next<= 23 ;
        245 : Address_next<= 46 ;
        247 : Address_next<= 47 ;
        248 : Address_next<= 23 ;
        249 : Address_next<= 11 ;
        250 : Address_next<= 5 ;
        251 : Address_next<= 2 ;
        254 : Address_next<= 3 ;
        255 : Address_next<= 6 ;
        256 : Address_next<= 12 ;
        257 : Address_next<= 24 ;
        258 : Address_next<= 48 ;
        260 : Address_next<= 49 ;
        261 : Address_next<= 24 ;
        263 : Address_next<= 25 ;
        264 : Address_next<= 50 ;
        266 : Address_next<= 51 ;
        267 : Address_next<= 25 ;
        268 : Address_next<= 12 ;
        270 : Address_next<= 13 ;
        271 : Address_next<= 26 ;
        272 : Address_next<= 52 ;
        274 : Address_next<= 53 ;
        275 : Address_next<= 26 ;
        277 : Address_next<= 27 ;
        278 : Address_next<= 54 ;
        280 : Address_next<= 55 ;
        281 : Address_next<= 27 ;
        282 : Address_next<= 13 ;
        283 : Address_next<= 6 ;
        285 : Address_next<= 7 ;
        286 : Address_next<= 14 ;
        287 : Address_next<= 28 ;
        288 : Address_next<= 56 ;
        290 : Address_next<= 57 ;
        291 : Address_next<= 28 ;
        293 : Address_next<= 29 ;
        294 : Address_next<= 58 ;
        296 : Address_next<= 59 ;
        297 : Address_next<= 29 ;
        298 : Address_next<= 14 ;
        300 : Address_next<= 15 ;
        301 : Address_next<= 30 ;
        302 : Address_next<= 60 ;
        304 : Address_next<= 61 ;
        305 : Address_next<= 30 ;
        307 : Address_next<= 31 ;
        308 : Address_next<= 62 ;
        310 : Address_next<= 63 ;
        311 : Address_next<= 31 ;
        312 : Address_next<= 15 ;
        313 : Address_next<= 7 ;
        314 : Address_next<= 3 ;
        315 : Address_next<= 1 ;
        316 : Address_next<= 1 ;
        329 : Address_next<= 1 ;
        330 : Address_next<= 1 ;
        331 : Address_next<= 1 ;
        332 : Address_next<= 1 ;
        333 : Address_next<= 2 ;
        334 : Address_next<= 2 ;
        335 : Address_next<= 4 ;
        336 : Address_next<= 8 ;
        337 : Address_next<= 16 ;
        338 : Address_next<= 32 ;
        339 : Address_next<= 64 ;
        341 : Address_next<= 65 ;
        342 : Address_next<= 32 ;
        344 : Address_next<= 33 ;
        345 : Address_next<= 66 ;
        347 : Address_next<= 67 ;
        348 : Address_next<= 33 ;
        349 : Address_next<= 16 ;
        351 : Address_next<= 17 ;
        352 : Address_next<= 34 ;
        353 : Address_next<= 68 ;
        355 : Address_next<= 69 ;
        356 : Address_next<= 34 ;
        358 : Address_next<= 35 ;
        359 : Address_next<= 70 ;
        361 : Address_next<= 71 ;
        362 : Address_next<= 35 ;
        363 : Address_next<= 17 ;
        364 : Address_next<= 8 ;
        366 : Address_next<= 9 ;
        367 : Address_next<= 18 ;
        368 : Address_next<= 36 ;
        369 : Address_next<= 72 ;
        371 : Address_next<= 73 ;
        372 : Address_next<= 36 ;
        374 : Address_next<= 37 ;
        375 : Address_next<= 74 ;
        377 : Address_next<= 75 ;
        378 : Address_next<= 37 ;
        379 : Address_next<= 18 ;
        381 : Address_next<= 19 ;
        382 : Address_next<= 38 ;
        383 : Address_next<= 76 ;
        385 : Address_next<= 77 ;
        386 : Address_next<= 38 ;
        388 : Address_next<= 39 ;
        389 : Address_next<= 78 ;
        391 : Address_next<= 79 ;
        392 : Address_next<= 39 ;
        393 : Address_next<= 19 ;
        394 : Address_next<= 9 ;
        395 : Address_next<= 4 ;
        398 : Address_next<= 5 ;
        399 : Address_next<= 10 ;
        400 : Address_next<= 20 ;
        401 : Address_next<= 40 ;
        402 : Address_next<= 80 ;
        404 : Address_next<= 81 ;
        405 : Address_next<= 40 ;
        407 : Address_next<= 41 ;
        408 : Address_next<= 82 ;
        410 : Address_next<= 83 ;
        411 : Address_next<= 41 ;
        412 : Address_next<= 20 ;
        414 : Address_next<= 21 ;
        415 : Address_next<= 42 ;
        416 : Address_next<= 84 ;
        418 : Address_next<= 85 ;
        419 : Address_next<= 42 ;
        421 : Address_next<= 43 ;
        422 : Address_next<= 86 ;
        424 : Address_next<= 87 ;
        425 : Address_next<= 43 ;
        426 : Address_next<= 21 ;
        427 : Address_next<= 10 ;
        429 : Address_next<= 11 ;
        430 : Address_next<= 22 ;
        431 : Address_next<= 44 ;
        432 : Address_next<= 88 ;
        434 : Address_next<= 89 ;
        435 : Address_next<= 44 ;
        437 : Address_next<= 45 ;
        438 : Address_next<= 90 ;
        440 : Address_next<= 91 ;
        441 : Address_next<= 45 ;
        442 : Address_next<= 22 ;
        444 : Address_next<= 23 ;
        445 : Address_next<= 46 ;
        446 : Address_next<= 92 ;
        448 : Address_next<= 93 ;
        449 : Address_next<= 46 ;
        451 : Address_next<= 47 ;
        452 : Address_next<= 94 ;
        454 : Address_next<= 95 ;
        455 : Address_next<= 47 ;
        456 : Address_next<= 23 ;
        457 : Address_next<= 11 ;
        458 : Address_next<= 5 ;
        459 : Address_next<= 2 ;
        460 : Address_next<= 2 ;
        465 : Address_next<= 3 ;
        466 : Address_next<= 3 ;
        467 : Address_next<= 6 ;
        468 : Address_next<= 12 ;
        469 : Address_next<= 24 ;
        470 : Address_next<= 48 ;
        471 : Address_next<= 96 ;
        473 : Address_next<= 97 ;
        474 : Address_next<= 48 ;
        476 : Address_next<= 49 ;
        477 : Address_next<= 98 ;
        479 : Address_next<= 99 ;
        480 : Address_next<= 49 ;
        481 : Address_next<= 24 ;
        483 : Address_next<= 25 ;
        484 : Address_next<= 50 ;
        485 : Address_next<= 100 ;
        487 : Address_next<= 101 ;
        488 : Address_next<= 50 ;
        490 : Address_next<= 51 ;
        491 : Address_next<= 102 ;
        493 : Address_next<= 103 ;
        494 : Address_next<= 51 ;
        495 : Address_next<= 25 ;
        496 : Address_next<= 12 ;
        498 : Address_next<= 13 ;
        499 : Address_next<= 26 ;
        500 : Address_next<= 52 ;
        501 : Address_next<= 104 ;
        503 : Address_next<= 105 ;
        504 : Address_next<= 52 ;
        506 : Address_next<= 53 ;
        507 : Address_next<= 106 ;
        509 : Address_next<= 107 ;
        510 : Address_next<= 53 ;
        511 : Address_next<= 26 ;
        513 : Address_next<= 27 ;
        514 : Address_next<= 54 ;
        515 : Address_next<= 108 ;
        517 : Address_next<= 109 ;
        518 : Address_next<= 54 ;
        520 : Address_next<= 55 ;
        521 : Address_next<= 110 ;
        523 : Address_next<= 111 ;
        524 : Address_next<= 55 ;
        525 : Address_next<= 27 ;
        526 : Address_next<= 13 ;
        527 : Address_next<= 6 ;
        530 : Address_next<= 7 ;
        531 : Address_next<= 14 ;
        532 : Address_next<= 28 ;
        533 : Address_next<= 56 ;
        534 : Address_next<= 112 ;
        536 : Address_next<= 113 ;
        537 : Address_next<= 56 ;
        539 : Address_next<= 57 ;
        540 : Address_next<= 114 ;
        542 : Address_next<= 115 ;
        543 : Address_next<= 57 ;
        544 : Address_next<= 28 ;
        546 : Address_next<= 29 ;
        547 : Address_next<= 58 ;
        548 : Address_next<= 116 ;
        550 : Address_next<= 117 ;
        551 : Address_next<= 58 ;
        553 : Address_next<= 59 ;
        554 : Address_next<= 118 ;
        556 : Address_next<= 119 ;
        557 : Address_next<= 59 ;
        558 : Address_next<= 29 ;
        559 : Address_next<= 14 ;
        561 : Address_next<= 15 ;
        562 : Address_next<= 30 ;
        563 : Address_next<= 60 ;
        564 : Address_next<= 120 ;
        566 : Address_next<= 121 ;
        567 : Address_next<= 60 ;
        569 : Address_next<= 61 ;
        570 : Address_next<= 122 ;
        572 : Address_next<= 123 ;
        573 : Address_next<= 61 ;
        574 : Address_next<= 30 ;
        576 : Address_next<= 31 ;
        577 : Address_next<= 62 ;
        578 : Address_next<= 124 ;
        580 : Address_next<= 125 ;
        581 : Address_next<= 62 ;
        583 : Address_next<= 63 ;
        584 : Address_next<= 126 ;
        586 : Address_next<= 127 ;
        587 : Address_next<= 63 ;
        588 : Address_next<= 31 ;
        589 : Address_next<= 15 ;
        590 : Address_next<= 7 ;
        591 : Address_next<= 3 ;
        592 : Address_next<= 3 ;
        593 : Address_next<= 1 ;
        594 : Address_next<= 1 ;
        595 : Address_next<= 1 ;
        596 : Address_next<= 1 ;
        621 : Address_next<= 1 ;
        622 : Address_next<= 1 ;
        623 : Address_next<= 1 ;
        624 : Address_next<= 1 ;
        625 : Address_next<= 1 ;
        626 : Address_next<= 1 ;
        627 : Address_next<= 1 ;
        628 : Address_next<= 1 ;
        629 : Address_next<= 2 ;
        630 : Address_next<= 2 ;
        631 : Address_next<= 2 ;
        632 : Address_next<= 2 ;
        633 : Address_next<= 4 ;
        634 : Address_next<= 4 ;
        635 : Address_next<= 8 ;
        636 : Address_next<= 16 ;
        637 : Address_next<= 32 ;
        638 : Address_next<= 64 ;
        639 : Address_next<= 128 ;
        641 : Address_next<= 129 ;
        642 : Address_next<= 64 ;
        644 : Address_next<= 65 ;
        645 : Address_next<= 130 ;
        647 : Address_next<= 131 ;
        648 : Address_next<= 65 ;
        649 : Address_next<= 32 ;
        651 : Address_next<= 33 ;
        652 : Address_next<= 66 ;
        653 : Address_next<= 132 ;
        655 : Address_next<= 133 ;
        656 : Address_next<= 66 ;
        658 : Address_next<= 67 ;
        659 : Address_next<= 134 ;
        661 : Address_next<= 135 ;
        662 : Address_next<= 67 ;
        663 : Address_next<= 33 ;
        664 : Address_next<= 16 ;
        666 : Address_next<= 17 ;
        667 : Address_next<= 34 ;
        668 : Address_next<= 68 ;
        669 : Address_next<= 136 ;
        671 : Address_next<= 137 ;
        672 : Address_next<= 68 ;
        674 : Address_next<= 69 ;
        675 : Address_next<= 138 ;
        677 : Address_next<= 139 ;
        678 : Address_next<= 69 ;
        679 : Address_next<= 34 ;
        681 : Address_next<= 35 ;
        682 : Address_next<= 70 ;
        683 : Address_next<= 140 ;
        685 : Address_next<= 141 ;
        686 : Address_next<= 70 ;
        688 : Address_next<= 71 ;
        689 : Address_next<= 142 ;
        691 : Address_next<= 143 ;
        692 : Address_next<= 71 ;
        693 : Address_next<= 35 ;
        694 : Address_next<= 17 ;
        695 : Address_next<= 8 ;
        698 : Address_next<= 9 ;
        699 : Address_next<= 18 ;
        700 : Address_next<= 36 ;
        701 : Address_next<= 72 ;
        702 : Address_next<= 144 ;
        704 : Address_next<= 145 ;
        705 : Address_next<= 72 ;
        707 : Address_next<= 73 ;
        708 : Address_next<= 146 ;
        710 : Address_next<= 147 ;
        711 : Address_next<= 73 ;
        712 : Address_next<= 36 ;
        714 : Address_next<= 37 ;
        715 : Address_next<= 74 ;
        716 : Address_next<= 148 ;
        718 : Address_next<= 149 ;
        719 : Address_next<= 74 ;
        721 : Address_next<= 75 ;
        722 : Address_next<= 150 ;
        724 : Address_next<= 151 ;
        725 : Address_next<= 75 ;
        726 : Address_next<= 37 ;
        727 : Address_next<= 18 ;
        729 : Address_next<= 19 ;
        730 : Address_next<= 38 ;
        731 : Address_next<= 76 ;
        732 : Address_next<= 152 ;
        734 : Address_next<= 153 ;
        735 : Address_next<= 76 ;
        737 : Address_next<= 77 ;
        738 : Address_next<= 154 ;
        740 : Address_next<= 155 ;
        741 : Address_next<= 77 ;
        742 : Address_next<= 38 ;
        744 : Address_next<= 39 ;
        745 : Address_next<= 78 ;
        746 : Address_next<= 156 ;
        748 : Address_next<= 157 ;
        749 : Address_next<= 78 ;
        751 : Address_next<= 79 ;
        752 : Address_next<= 158 ;
        754 : Address_next<= 159 ;
        755 : Address_next<= 79 ;
        756 : Address_next<= 39 ;
        757 : Address_next<= 19 ;
        758 : Address_next<= 9 ;
        759 : Address_next<= 4 ;
        760 : Address_next<= 4 ;
        765 : Address_next<= 5 ;
        766 : Address_next<= 5 ;
        767 : Address_next<= 10 ;
        768 : Address_next<= 20 ;
        769 : Address_next<= 40 ;
        770 : Address_next<= 80 ;
        771 : Address_next<= 160 ;
        773 : Address_next<= 161 ;
        774 : Address_next<= 80 ;
        776 : Address_next<= 81 ;
        777 : Address_next<= 162 ;
        779 : Address_next<= 163 ;
        780 : Address_next<= 81 ;
        781 : Address_next<= 40 ;
        783 : Address_next<= 41 ;
        784 : Address_next<= 82 ;
        785 : Address_next<= 164 ;
        787 : Address_next<= 165 ;
        788 : Address_next<= 82 ;
        790 : Address_next<= 83 ;
        791 : Address_next<= 166 ;
        793 : Address_next<= 167 ;
        794 : Address_next<= 83 ;
        795 : Address_next<= 41 ;
        796 : Address_next<= 20 ;
        798 : Address_next<= 21 ;
        799 : Address_next<= 42 ;
        800 : Address_next<= 84 ;
        801 : Address_next<= 168 ;
        803 : Address_next<= 169 ;
        804 : Address_next<= 84 ;
        806 : Address_next<= 85 ;
        807 : Address_next<= 170 ;
        809 : Address_next<= 171 ;
        810 : Address_next<= 85 ;
        811 : Address_next<= 42 ;
        813 : Address_next<= 43 ;
        814 : Address_next<= 86 ;
        815 : Address_next<= 172 ;
        817 : Address_next<= 173 ;
        818 : Address_next<= 86 ;
        820 : Address_next<= 87 ;
        821 : Address_next<= 174 ;
        823 : Address_next<= 175 ;
        824 : Address_next<= 87 ;
        825 : Address_next<= 43 ;
        826 : Address_next<= 21 ;
        827 : Address_next<= 10 ;
        830 : Address_next<= 11 ;
        831 : Address_next<= 22 ;
        832 : Address_next<= 44 ;
        833 : Address_next<= 88 ;
        834 : Address_next<= 176 ;
        836 : Address_next<= 177 ;
        837 : Address_next<= 88 ;
        839 : Address_next<= 89 ;
        840 : Address_next<= 178 ;
        842 : Address_next<= 179 ;
        843 : Address_next<= 89 ;
        844 : Address_next<= 44 ;
        846 : Address_next<= 45 ;
        847 : Address_next<= 90 ;
        848 : Address_next<= 180 ;
        850 : Address_next<= 181 ;
        851 : Address_next<= 90 ;
        853 : Address_next<= 91 ;
        854 : Address_next<= 182 ;
        856 : Address_next<= 183 ;
        857 : Address_next<= 91 ;
        858 : Address_next<= 45 ;
        859 : Address_next<= 22 ;
        861 : Address_next<= 23 ;
        862 : Address_next<= 46 ;
        863 : Address_next<= 92 ;
        864 : Address_next<= 184 ;
        866 : Address_next<= 185 ;
        867 : Address_next<= 92 ;
        869 : Address_next<= 93 ;
        870 : Address_next<= 186 ;
        872 : Address_next<= 187 ;
        873 : Address_next<= 93 ;
        874 : Address_next<= 46 ;
        876 : Address_next<= 47 ;
        877 : Address_next<= 94 ;
        878 : Address_next<= 188 ;
        880 : Address_next<= 189 ;
        881 : Address_next<= 94 ;
        883 : Address_next<= 95 ;
        884 : Address_next<= 190 ;
        886 : Address_next<= 191 ;
        887 : Address_next<= 95 ;
        888 : Address_next<= 47 ;
        889 : Address_next<= 23 ;
        890 : Address_next<= 11 ;
        891 : Address_next<= 5 ;
        892 : Address_next<= 5 ;
        893 : Address_next<= 2 ;
        894 : Address_next<= 2 ;
        895 : Address_next<= 2 ;
        896 : Address_next<= 2 ;
        905 : Address_next<= 3 ;
        906 : Address_next<= 3 ;
        907 : Address_next<= 3 ;
        908 : Address_next<= 3 ;
        909 : Address_next<= 6 ;
        910 : Address_next<= 6 ;
        911 : Address_next<= 12 ;
        912 : Address_next<= 24 ;
        913 : Address_next<= 48 ;
        914 : Address_next<= 96 ;
        915 : Address_next<= 192 ;
        917 : Address_next<= 193 ;
        918 : Address_next<= 96 ;
        920 : Address_next<= 97 ;
        921 : Address_next<= 194 ;
        923 : Address_next<= 195 ;
        924 : Address_next<= 97 ;
        925 : Address_next<= 48 ;
        927 : Address_next<= 49 ;
        928 : Address_next<= 98 ;
        929 : Address_next<= 196 ;
        931 : Address_next<= 197 ;
        932 : Address_next<= 98 ;
        934 : Address_next<= 99 ;
        935 : Address_next<= 198 ;
        937 : Address_next<= 199 ;
        938 : Address_next<= 99 ;
        939 : Address_next<= 49 ;
        940 : Address_next<= 24 ;
        942 : Address_next<= 25 ;
        943 : Address_next<= 50 ;
        944 : Address_next<= 100 ;
        945 : Address_next<= 200 ;
        947 : Address_next<= 201 ;
        948 : Address_next<= 100 ;
        950 : Address_next<= 101 ;
        951 : Address_next<= 202 ;
        953 : Address_next<= 203 ;
        954 : Address_next<= 101 ;
        955 : Address_next<= 50 ;
        957 : Address_next<= 51 ;
        958 : Address_next<= 102 ;
        959 : Address_next<= 204 ;
        961 : Address_next<= 205 ;
        962 : Address_next<= 102 ;
        964 : Address_next<= 103 ;
        965 : Address_next<= 206 ;
        967 : Address_next<= 207 ;
        968 : Address_next<= 103 ;
        969 : Address_next<= 51 ;
        970 : Address_next<= 25 ;
        971 : Address_next<= 12 ;
        974 : Address_next<= 13 ;
        975 : Address_next<= 26 ;
        976 : Address_next<= 52 ;
        977 : Address_next<= 104 ;
        978 : Address_next<= 208 ;
        980 : Address_next<= 209 ;
        981 : Address_next<= 104 ;
        983 : Address_next<= 105 ;
        984 : Address_next<= 210 ;
        986 : Address_next<= 211 ;
        987 : Address_next<= 105 ;
        988 : Address_next<= 52 ;
        990 : Address_next<= 53 ;
        991 : Address_next<= 106 ;
        992 : Address_next<= 212 ;
        994 : Address_next<= 213 ;
        995 : Address_next<= 106 ;
        997 : Address_next<= 107 ;
        998 : Address_next<= 214 ;
        1000 : Address_next<= 215 ;
        1001 : Address_next<= 107 ;
        1002 : Address_next<= 53 ;
        1003 : Address_next<= 26 ;
        1005 : Address_next<= 27 ;
        1006 : Address_next<= 54 ;
        1007 : Address_next<= 108 ;
        1008 : Address_next<= 216 ;
        1010 : Address_next<= 217 ;
        1011 : Address_next<= 108 ;
        1013 : Address_next<= 109 ;
        1014 : Address_next<= 218 ;
        1016 : Address_next<= 219 ;
        1017 : Address_next<= 109 ;
        1018 : Address_next<= 54 ;
        1020 : Address_next<= 55 ;
        1021 : Address_next<= 110 ;
        1022 : Address_next<= 220 ;
        1024 : Address_next<= 221 ;
        1025 : Address_next<= 110 ;
        1027 : Address_next<= 111 ;
        1028 : Address_next<= 222 ;
        1030 : Address_next<= 223 ;
        1031 : Address_next<= 111 ;
        1032 : Address_next<= 55 ;
        1033 : Address_next<= 27 ;
        1034 : Address_next<= 13 ;
        1035 : Address_next<= 6 ;
        1036 : Address_next<= 6 ;
        1041 : Address_next<= 7 ;
        1042 : Address_next<= 7 ;
        1043 : Address_next<= 14 ;
        1044 : Address_next<= 28 ;
        1045 : Address_next<= 56 ;
        1046 : Address_next<= 112 ;
        1047 : Address_next<= 224 ;
        1049 : Address_next<= 225 ;
        1050 : Address_next<= 112 ;
        1052 : Address_next<= 113 ;
        1053 : Address_next<= 226 ;
        1055 : Address_next<= 227 ;
        1056 : Address_next<= 113 ;
        1057 : Address_next<= 56 ;
        1059 : Address_next<= 57 ;
        1060 : Address_next<= 114 ;
        1061 : Address_next<= 228 ;
        1063 : Address_next<= 229 ;
        1064 : Address_next<= 114 ;
        1066 : Address_next<= 115 ;
        1067 : Address_next<= 230 ;
        1069 : Address_next<= 231 ;
        1070 : Address_next<= 115 ;
        1071 : Address_next<= 57 ;
        1072 : Address_next<= 28 ;
        1074 : Address_next<= 29 ;
        1075 : Address_next<= 58 ;
        1076 : Address_next<= 116 ;
        1077 : Address_next<= 232 ;
        1079 : Address_next<= 233 ;
        1080 : Address_next<= 116 ;
        1082 : Address_next<= 117 ;
        1083 : Address_next<= 234 ;
        1085 : Address_next<= 235 ;
        1086 : Address_next<= 117 ;
        1087 : Address_next<= 58 ;
        1089 : Address_next<= 59 ;
        1090 : Address_next<= 118 ;
        1091 : Address_next<= 236 ;
        1093 : Address_next<= 237 ;
        1094 : Address_next<= 118 ;
        1096 : Address_next<= 119 ;
        1097 : Address_next<= 238 ;
        1099 : Address_next<= 239 ;
        1100 : Address_next<= 119 ;
        1101 : Address_next<= 59 ;
        1102 : Address_next<= 29 ;
        1103 : Address_next<= 14 ;
        1106 : Address_next<= 15 ;
        1107 : Address_next<= 30 ;
        1108 : Address_next<= 60 ;
        1109 : Address_next<= 120 ;
        1110 : Address_next<= 240 ;
        1112 : Address_next<= 241 ;
        1113 : Address_next<= 120 ;
        1115 : Address_next<= 121 ;
        1116 : Address_next<= 242 ;
        1118 : Address_next<= 243 ;
        1119 : Address_next<= 121 ;
        1120 : Address_next<= 60 ;
        1122 : Address_next<= 61 ;
        1123 : Address_next<= 122 ;
        1124 : Address_next<= 244 ;
        1126 : Address_next<= 245 ;
        1127 : Address_next<= 122 ;
        1129 : Address_next<= 123 ;
        1130 : Address_next<= 246 ;
        1132 : Address_next<= 247 ;
        1133 : Address_next<= 123 ;
        1134 : Address_next<= 61 ;
        1135 : Address_next<= 30 ;
        1137 : Address_next<= 31 ;
        1138 : Address_next<= 62 ;
        1139 : Address_next<= 124 ;
        1140 : Address_next<= 248 ;
        1142 : Address_next<= 249 ;
        1143 : Address_next<= 124 ;
        1145 : Address_next<= 125 ;
        1146 : Address_next<= 250 ;
        1148 : Address_next<= 251 ;
        1149 : Address_next<= 125 ;
        1150 : Address_next<= 62 ;
        1152 : Address_next<= 63 ;
        1153 : Address_next<= 126 ;
        1154 : Address_next<= 252 ;
        1156 : Address_next<= 253 ;
        1157 : Address_next<= 126 ;
        1159 : Address_next<= 127 ;
        1160 : Address_next<= 254 ;
        1162 : Address_next<= 255 ;
        1163 : Address_next<= 127 ;
        1164 : Address_next<= 63 ;
        1165 : Address_next<= 31 ;
        1166 : Address_next<= 15 ;
        1167 : Address_next<= 7 ;
        1168 : Address_next<= 7 ;
        1169 : Address_next<= 3 ;
        1170 : Address_next<= 3 ;
        1171 : Address_next<= 3 ;
        1172 : Address_next<= 3 ;
        1173 : Address_next<= 1 ;
        1174 : Address_next<= 1 ;
        1175 : Address_next<= 1 ;
        1176 : Address_next<= 1 ;
        1177 : Address_next<= 1 ;
        1178 : Address_next<= 1 ;
        1179 : Address_next<= 1 ;
        1180 : Address_next<= 1 ;
        1229 : Address_next<= 1 ;
        1230 : Address_next<= 1 ;
        1231 : Address_next<= 1 ;
        1232 : Address_next<= 1 ;
        1233 : Address_next<= 1 ;
        1234 : Address_next<= 1 ;
        1235 : Address_next<= 1 ;
        1236 : Address_next<= 1 ;
        1237 : Address_next<= 1 ;
        1238 : Address_next<= 1 ;
        1239 : Address_next<= 1 ;
        1240 : Address_next<= 1 ;
        1241 : Address_next<= 1 ;
        1242 : Address_next<= 1 ;
        1243 : Address_next<= 1 ;
        1244 : Address_next<= 1 ;
        1245 : Address_next<= 2 ;
        1246 : Address_next<= 2 ;
        1247 : Address_next<= 2 ;
        1248 : Address_next<= 2 ;
        1249 : Address_next<= 2 ;
        1250 : Address_next<= 2 ;
        1251 : Address_next<= 2 ;
        1252 : Address_next<= 2 ;
        1253 : Address_next<= 4 ;
        1254 : Address_next<= 4 ;
        1255 : Address_next<= 4 ;
        1256 : Address_next<= 4 ;
        1257 : Address_next<= 8 ;
        1258 : Address_next<= 8 ;
        1259 : Address_next<= 16 ;
        1260 : Address_next<= 32 ;
        1261 : Address_next<= 64 ;
        1262 : Address_next<= 128 ;
        1263 : Address_next<= 256 ;
        1265 : Address_next<= 257 ;
        1266 : Address_next<= 128 ;
        1268 : Address_next<= 129 ;
        1269 : Address_next<= 258 ;
        1271 : Address_next<= 259 ;
        1272 : Address_next<= 129 ;
        1273 : Address_next<= 64 ;
        1275 : Address_next<= 65 ;
        1276 : Address_next<= 130 ;
        1277 : Address_next<= 260 ;
        1279 : Address_next<= 261 ;
        1280 : Address_next<= 130 ;
        1282 : Address_next<= 131 ;
        1283 : Address_next<= 262 ;
        1285 : Address_next<= 263 ;
        1286 : Address_next<= 131 ;
        1287 : Address_next<= 65 ;
        1288 : Address_next<= 32 ;
        1290 : Address_next<= 33 ;
        1291 : Address_next<= 66 ;
        1292 : Address_next<= 132 ;
        1293 : Address_next<= 264 ;
        1295 : Address_next<= 265 ;
        1296 : Address_next<= 132 ;
        1298 : Address_next<= 133 ;
        1299 : Address_next<= 266 ;
        1301 : Address_next<= 267 ;
        1302 : Address_next<= 133 ;
        1303 : Address_next<= 66 ;
        1305 : Address_next<= 67 ;
        1306 : Address_next<= 134 ;
        1307 : Address_next<= 268 ;
        1309 : Address_next<= 269 ;
        1310 : Address_next<= 134 ;
        1312 : Address_next<= 135 ;
        1313 : Address_next<= 270 ;
        1315 : Address_next<= 271 ;
        1316 : Address_next<= 135 ;
        1317 : Address_next<= 67 ;
        1318 : Address_next<= 33 ;
        1319 : Address_next<= 16 ;
        1322 : Address_next<= 17 ;
        1323 : Address_next<= 34 ;
        1324 : Address_next<= 68 ;
        1325 : Address_next<= 136 ;
        1326 : Address_next<= 272 ;
        1328 : Address_next<= 273 ;
        1329 : Address_next<= 136 ;
        1331 : Address_next<= 137 ;
        1332 : Address_next<= 274 ;
        1334 : Address_next<= 275 ;
        1335 : Address_next<= 137 ;
        1336 : Address_next<= 68 ;
        1338 : Address_next<= 69 ;
        1339 : Address_next<= 138 ;
        1340 : Address_next<= 276 ;
        1342 : Address_next<= 277 ;
        1343 : Address_next<= 138 ;
        1345 : Address_next<= 139 ;
        1346 : Address_next<= 278 ;
        1348 : Address_next<= 279 ;
        1349 : Address_next<= 139 ;
        1350 : Address_next<= 69 ;
        1351 : Address_next<= 34 ;
        1353 : Address_next<= 35 ;
        1354 : Address_next<= 70 ;
        1355 : Address_next<= 140 ;
        1356 : Address_next<= 280 ;
        1358 : Address_next<= 281 ;
        1359 : Address_next<= 140 ;
        1361 : Address_next<= 141 ;
        1362 : Address_next<= 282 ;
        1364 : Address_next<= 283 ;
        1365 : Address_next<= 141 ;
        1366 : Address_next<= 70 ;
        1368 : Address_next<= 71 ;
        1369 : Address_next<= 142 ;
        1370 : Address_next<= 284 ;
        1372 : Address_next<= 285 ;
        1373 : Address_next<= 142 ;
        1375 : Address_next<= 143 ;
        1376 : Address_next<= 286 ;
        1378 : Address_next<= 287 ;
        1379 : Address_next<= 143 ;
        1380 : Address_next<= 71 ;
        1381 : Address_next<= 35 ;
        1382 : Address_next<= 17 ;
        1383 : Address_next<= 8 ;
        1384 : Address_next<= 8 ;
        1389 : Address_next<= 9 ;
        1390 : Address_next<= 9 ;
        1391 : Address_next<= 18 ;
        1392 : Address_next<= 36 ;
        1393 : Address_next<= 72 ;
        1394 : Address_next<= 144 ;
        1395 : Address_next<= 288 ;
        1397 : Address_next<= 289 ;
        1398 : Address_next<= 144 ;
        1400 : Address_next<= 145 ;
        1401 : Address_next<= 290 ;
        1403 : Address_next<= 291 ;
        1404 : Address_next<= 145 ;
        1405 : Address_next<= 72 ;
        1407 : Address_next<= 73 ;
        1408 : Address_next<= 146 ;
        1409 : Address_next<= 292 ;
        1411 : Address_next<= 293 ;
        1412 : Address_next<= 146 ;
        1414 : Address_next<= 147 ;
        1415 : Address_next<= 294 ;
        1417 : Address_next<= 295 ;
        1418 : Address_next<= 147 ;
        1419 : Address_next<= 73 ;
        1420 : Address_next<= 36 ;
        1422 : Address_next<= 37 ;
        1423 : Address_next<= 74 ;
        1424 : Address_next<= 148 ;
        1425 : Address_next<= 296 ;
        1427 : Address_next<= 297 ;
        1428 : Address_next<= 148 ;
        1430 : Address_next<= 149 ;
        1431 : Address_next<= 298 ;
        1433 : Address_next<= 299 ;
        1434 : Address_next<= 149 ;
        1435 : Address_next<= 74 ;
        1437 : Address_next<= 75 ;
        1438 : Address_next<= 150 ;
        1439 : Address_next<= 300 ;
        1441 : Address_next<= 301 ;
        1442 : Address_next<= 150 ;
        1444 : Address_next<= 151 ;
        1445 : Address_next<= 302 ;
        1447 : Address_next<= 303 ;
        1448 : Address_next<= 151 ;
        1449 : Address_next<= 75 ;
        1450 : Address_next<= 37 ;
        1451 : Address_next<= 18 ;
        1454 : Address_next<= 19 ;
        1455 : Address_next<= 38 ;
        1456 : Address_next<= 76 ;
        1457 : Address_next<= 152 ;
        1458 : Address_next<= 304 ;
        1460 : Address_next<= 305 ;
        1461 : Address_next<= 152 ;
        1463 : Address_next<= 153 ;
        1464 : Address_next<= 306 ;
        1466 : Address_next<= 307 ;
        1467 : Address_next<= 153 ;
        1468 : Address_next<= 76 ;
        1470 : Address_next<= 77 ;
        1471 : Address_next<= 154 ;
        1472 : Address_next<= 308 ;
        1474 : Address_next<= 309 ;
        1475 : Address_next<= 154 ;
        1477 : Address_next<= 155 ;
        1478 : Address_next<= 310 ;
        1480 : Address_next<= 311 ;
        1481 : Address_next<= 155 ;
        1482 : Address_next<= 77 ;
        1483 : Address_next<= 38 ;
        1485 : Address_next<= 39 ;
        1486 : Address_next<= 78 ;
        1487 : Address_next<= 156 ;
        1488 : Address_next<= 312 ;
        1490 : Address_next<= 313 ;
        1491 : Address_next<= 156 ;
        1493 : Address_next<= 157 ;
        1494 : Address_next<= 314 ;
        1496 : Address_next<= 315 ;
        1497 : Address_next<= 157 ;
        1498 : Address_next<= 78 ;
        1500 : Address_next<= 79 ;
        1501 : Address_next<= 158 ;
        1502 : Address_next<= 316 ;
        1504 : Address_next<= 317 ;
        1505 : Address_next<= 158 ;
        1507 : Address_next<= 159 ;
        1508 : Address_next<= 318 ;
        1510 : Address_next<= 319 ;
        1511 : Address_next<= 159 ;
        1512 : Address_next<= 79 ;
        1513 : Address_next<= 39 ;
        1514 : Address_next<= 19 ;
        1515 : Address_next<= 9 ;
        1516 : Address_next<= 9 ;
        1517 : Address_next<= 4 ;
        1518 : Address_next<= 4 ;
        1519 : Address_next<= 4 ;
        1520 : Address_next<= 4 ;
        1529 : Address_next<= 5 ;
        1530 : Address_next<= 5 ;
        1531 : Address_next<= 5 ;
        1532 : Address_next<= 5 ;
        1533 : Address_next<= 10 ;
        1534 : Address_next<= 10 ;
        1535 : Address_next<= 20 ;
        1536 : Address_next<= 40 ;
        1537 : Address_next<= 80 ;
        1538 : Address_next<= 160 ;
        1539 : Address_next<= 320 ;
        1541 : Address_next<= 321 ;
        1542 : Address_next<= 160 ;
        1544 : Address_next<= 161 ;
        1545 : Address_next<= 322 ;
        1547 : Address_next<= 323 ;
        1548 : Address_next<= 161 ;
        1549 : Address_next<= 80 ;
        1551 : Address_next<= 81 ;
        1552 : Address_next<= 162 ;
        1553 : Address_next<= 324 ;
        1555 : Address_next<= 325 ;
        1556 : Address_next<= 162 ;
        1558 : Address_next<= 163 ;
        1559 : Address_next<= 326 ;
        1561 : Address_next<= 327 ;
        1562 : Address_next<= 163 ;
        1563 : Address_next<= 81 ;
        1564 : Address_next<= 40 ;
        1566 : Address_next<= 41 ;
        1567 : Address_next<= 82 ;
        1568 : Address_next<= 164 ;
        1569 : Address_next<= 328 ;
        1571 : Address_next<= 329 ;
        1572 : Address_next<= 164 ;
        1574 : Address_next<= 165 ;
        1575 : Address_next<= 330 ;
        1577 : Address_next<= 331 ;
        1578 : Address_next<= 165 ;
        1579 : Address_next<= 82 ;
        1581 : Address_next<= 83 ;
        1582 : Address_next<= 166 ;
        1583 : Address_next<= 332 ;
        1585 : Address_next<= 333 ;
        1586 : Address_next<= 166 ;
        1588 : Address_next<= 167 ;
        1589 : Address_next<= 334 ;
        1591 : Address_next<= 335 ;
        1592 : Address_next<= 167 ;
        1593 : Address_next<= 83 ;
        1594 : Address_next<= 41 ;
        1595 : Address_next<= 20 ;
        1598 : Address_next<= 21 ;
        1599 : Address_next<= 42 ;
        1600 : Address_next<= 84 ;
        1601 : Address_next<= 168 ;
        1602 : Address_next<= 336 ;
        1604 : Address_next<= 337 ;
        1605 : Address_next<= 168 ;
        1607 : Address_next<= 169 ;
        1608 : Address_next<= 338 ;
        1610 : Address_next<= 339 ;
        1611 : Address_next<= 169 ;
        1612 : Address_next<= 84 ;
        1614 : Address_next<= 85 ;
        1615 : Address_next<= 170 ;
        1616 : Address_next<= 340 ;
        1618 : Address_next<= 341 ;
        1619 : Address_next<= 170 ;
        1621 : Address_next<= 171 ;
        1622 : Address_next<= 342 ;
        1624 : Address_next<= 343 ;
        1625 : Address_next<= 171 ;
        1626 : Address_next<= 85 ;
        1627 : Address_next<= 42 ;
        1629 : Address_next<= 43 ;
        1630 : Address_next<= 86 ;
        1631 : Address_next<= 172 ;
        1632 : Address_next<= 344 ;
        1634 : Address_next<= 345 ;
        1635 : Address_next<= 172 ;
        1637 : Address_next<= 173 ;
        1638 : Address_next<= 346 ;
        1640 : Address_next<= 347 ;
        1641 : Address_next<= 173 ;
        1642 : Address_next<= 86 ;
        1644 : Address_next<= 87 ;
        1645 : Address_next<= 174 ;
        1646 : Address_next<= 348 ;
        1648 : Address_next<= 349 ;
        1649 : Address_next<= 174 ;
        1651 : Address_next<= 175 ;
        1652 : Address_next<= 350 ;
        1654 : Address_next<= 351 ;
        1655 : Address_next<= 175 ;
        1656 : Address_next<= 87 ;
        1657 : Address_next<= 43 ;
        1658 : Address_next<= 21 ;
        1659 : Address_next<= 10 ;
        1660 : Address_next<= 10 ;
        1665 : Address_next<= 11 ;
        1666 : Address_next<= 11 ;
        1667 : Address_next<= 22 ;
        1668 : Address_next<= 44 ;
        1669 : Address_next<= 88 ;
        1670 : Address_next<= 176 ;
        1671 : Address_next<= 352 ;
        1673 : Address_next<= 353 ;
        1674 : Address_next<= 176 ;
        1676 : Address_next<= 177 ;
        1677 : Address_next<= 354 ;
        1679 : Address_next<= 355 ;
        1680 : Address_next<= 177 ;
        1681 : Address_next<= 88 ;
        1683 : Address_next<= 89 ;
        1684 : Address_next<= 178 ;
        1685 : Address_next<= 356 ;
        1687 : Address_next<= 357 ;
        1688 : Address_next<= 178 ;
        1690 : Address_next<= 179 ;
        1691 : Address_next<= 358 ;
        1693 : Address_next<= 359 ;
        1694 : Address_next<= 179 ;
        1695 : Address_next<= 89 ;
        1696 : Address_next<= 44 ;
        1698 : Address_next<= 45 ;
        1699 : Address_next<= 90 ;
        1700 : Address_next<= 180 ;
        1701 : Address_next<= 360 ;
        1703 : Address_next<= 361 ;
        1704 : Address_next<= 180 ;
        1706 : Address_next<= 181 ;
        1707 : Address_next<= 362 ;
        1709 : Address_next<= 363 ;
        1710 : Address_next<= 181 ;
        1711 : Address_next<= 90 ;
        1713 : Address_next<= 91 ;
        1714 : Address_next<= 182 ;
        1715 : Address_next<= 364 ;
        1717 : Address_next<= 365 ;
        1718 : Address_next<= 182 ;
        1720 : Address_next<= 183 ;
        1721 : Address_next<= 366 ;
        1723 : Address_next<= 367 ;
        1724 : Address_next<= 183 ;
        1725 : Address_next<= 91 ;
        1726 : Address_next<= 45 ;
        1727 : Address_next<= 22 ;
        1730 : Address_next<= 23 ;
        1731 : Address_next<= 46 ;
        1732 : Address_next<= 92 ;
        1733 : Address_next<= 184 ;
        1734 : Address_next<= 368 ;
        1736 : Address_next<= 369 ;
        1737 : Address_next<= 184 ;
        1739 : Address_next<= 185 ;
        1740 : Address_next<= 370 ;
        1742 : Address_next<= 371 ;
        1743 : Address_next<= 185 ;
        1744 : Address_next<= 92 ;
        1746 : Address_next<= 93 ;
        1747 : Address_next<= 186 ;
        1748 : Address_next<= 372 ;
        1750 : Address_next<= 373 ;
        1751 : Address_next<= 186 ;
        1753 : Address_next<= 187 ;
        1754 : Address_next<= 374 ;
        1756 : Address_next<= 375 ;
        1757 : Address_next<= 187 ;
        1758 : Address_next<= 93 ;
        1759 : Address_next<= 46 ;
        1761 : Address_next<= 47 ;
        1762 : Address_next<= 94 ;
        1763 : Address_next<= 188 ;
        1764 : Address_next<= 376 ;
        1766 : Address_next<= 377 ;
        1767 : Address_next<= 188 ;
        1769 : Address_next<= 189 ;
        1770 : Address_next<= 378 ;
        1772 : Address_next<= 379 ;
        1773 : Address_next<= 189 ;
        1774 : Address_next<= 94 ;
        1776 : Address_next<= 95 ;
        1777 : Address_next<= 190 ;
        1778 : Address_next<= 380 ;
        1780 : Address_next<= 381 ;
        1781 : Address_next<= 190 ;
        1783 : Address_next<= 191 ;
        1784 : Address_next<= 382 ;
        1786 : Address_next<= 383 ;
        1787 : Address_next<= 191 ;
        1788 : Address_next<= 95 ;
        1789 : Address_next<= 47 ;
        1790 : Address_next<= 23 ;
        1791 : Address_next<= 11 ;
        1792 : Address_next<= 11 ;
        1793 : Address_next<= 5 ;
        1794 : Address_next<= 5 ;
        1795 : Address_next<= 5 ;
        1796 : Address_next<= 5 ;
        1797 : Address_next<= 2 ;
        1798 : Address_next<= 2 ;
        1799 : Address_next<= 2 ;
        1800 : Address_next<= 2 ;
        1801 : Address_next<= 2 ;
        1802 : Address_next<= 2 ;
        1803 : Address_next<= 2 ;
        1804 : Address_next<= 2 ;
        1821 : Address_next<= 3 ;
        1822 : Address_next<= 3 ;
        1823 : Address_next<= 3 ;
        1824 : Address_next<= 3 ;
        1825 : Address_next<= 3 ;
        1826 : Address_next<= 3 ;
        1827 : Address_next<= 3 ;
        1828 : Address_next<= 3 ;
        1829 : Address_next<= 6 ;
        1830 : Address_next<= 6 ;
        1831 : Address_next<= 6 ;
        1832 : Address_next<= 6 ;
        1833 : Address_next<= 12 ;
        1834 : Address_next<= 12 ;
        1835 : Address_next<= 24 ;
        1836 : Address_next<= 48 ;
        1837 : Address_next<= 96 ;
        1838 : Address_next<= 192 ;
        1839 : Address_next<= 384 ;
        1841 : Address_next<= 385 ;
        1842 : Address_next<= 192 ;
        1844 : Address_next<= 193 ;
        1845 : Address_next<= 386 ;
        1847 : Address_next<= 387 ;
        1848 : Address_next<= 193 ;
        1849 : Address_next<= 96 ;
        1851 : Address_next<= 97 ;
        1852 : Address_next<= 194 ;
        1853 : Address_next<= 388 ;
        1855 : Address_next<= 389 ;
        1856 : Address_next<= 194 ;
        1858 : Address_next<= 195 ;
        1859 : Address_next<= 390 ;
        1861 : Address_next<= 391 ;
        1862 : Address_next<= 195 ;
        1863 : Address_next<= 97 ;
        1864 : Address_next<= 48 ;
        1866 : Address_next<= 49 ;
        1867 : Address_next<= 98 ;
        1868 : Address_next<= 196 ;
        1869 : Address_next<= 392 ;
        1871 : Address_next<= 393 ;
        1872 : Address_next<= 196 ;
        1874 : Address_next<= 197 ;
        1875 : Address_next<= 394 ;
        1877 : Address_next<= 395 ;
        1878 : Address_next<= 197 ;
        1879 : Address_next<= 98 ;
        1881 : Address_next<= 99 ;
        1882 : Address_next<= 198 ;
        1883 : Address_next<= 396 ;
        1885 : Address_next<= 397 ;
        1886 : Address_next<= 198 ;
        1888 : Address_next<= 199 ;
        1889 : Address_next<= 398 ;
        1891 : Address_next<= 399 ;
        1892 : Address_next<= 199 ;
        1893 : Address_next<= 99 ;
        1894 : Address_next<= 49 ;
        1895 : Address_next<= 24 ;
        1898 : Address_next<= 25 ;
        1899 : Address_next<= 50 ;
        1900 : Address_next<= 100 ;
        1901 : Address_next<= 200 ;
        1902 : Address_next<= 400 ;
        1904 : Address_next<= 401 ;
        1905 : Address_next<= 200 ;
        1907 : Address_next<= 201 ;
        1908 : Address_next<= 402 ;
        1910 : Address_next<= 403 ;
        1911 : Address_next<= 201 ;
        1912 : Address_next<= 100 ;
        1914 : Address_next<= 101 ;
        1915 : Address_next<= 202 ;
        1916 : Address_next<= 404 ;
        1918 : Address_next<= 405 ;
        1919 : Address_next<= 202 ;
        1921 : Address_next<= 203 ;
        1922 : Address_next<= 406 ;
        1924 : Address_next<= 407 ;
        1925 : Address_next<= 203 ;
        1926 : Address_next<= 101 ;
        1927 : Address_next<= 50 ;
        1929 : Address_next<= 51 ;
        1930 : Address_next<= 102 ;
        1931 : Address_next<= 204 ;
        1932 : Address_next<= 408 ;
        1934 : Address_next<= 409 ;
        1935 : Address_next<= 204 ;
        1937 : Address_next<= 205 ;
        1938 : Address_next<= 410 ;
        1940 : Address_next<= 411 ;
        1941 : Address_next<= 205 ;
        1942 : Address_next<= 102 ;
        1944 : Address_next<= 103 ;
        1945 : Address_next<= 206 ;
        1946 : Address_next<= 412 ;
        1948 : Address_next<= 413 ;
        1949 : Address_next<= 206 ;
        1951 : Address_next<= 207 ;
        1952 : Address_next<= 414 ;
        1954 : Address_next<= 415 ;
        1955 : Address_next<= 207 ;
        1956 : Address_next<= 103 ;
        1957 : Address_next<= 51 ;
        1958 : Address_next<= 25 ;
        1959 : Address_next<= 12 ;
        1960 : Address_next<= 12 ;
        1965 : Address_next<= 13 ;
        1966 : Address_next<= 13 ;
        1967 : Address_next<= 26 ;
        1968 : Address_next<= 52 ;
        1969 : Address_next<= 104 ;
        1970 : Address_next<= 208 ;
        1971 : Address_next<= 416 ;
        1973 : Address_next<= 417 ;
        1974 : Address_next<= 208 ;
        1976 : Address_next<= 209 ;
        1977 : Address_next<= 418 ;
        1979 : Address_next<= 419 ;
        1980 : Address_next<= 209 ;
        1981 : Address_next<= 104 ;
        1983 : Address_next<= 105 ;
        1984 : Address_next<= 210 ;
        1985 : Address_next<= 420 ;
        1987 : Address_next<= 421 ;
        1988 : Address_next<= 210 ;
        1990 : Address_next<= 211 ;
        1991 : Address_next<= 422 ;
        1993 : Address_next<= 423 ;
        1994 : Address_next<= 211 ;
        1995 : Address_next<= 105 ;
        1996 : Address_next<= 52 ;
        1998 : Address_next<= 53 ;
        1999 : Address_next<= 106 ;
        2000 : Address_next<= 212 ;
        2001 : Address_next<= 424 ;
        2003 : Address_next<= 425 ;
        2004 : Address_next<= 212 ;
        2006 : Address_next<= 213 ;
        2007 : Address_next<= 426 ;
        2009 : Address_next<= 427 ;
        2010 : Address_next<= 213 ;
        2011 : Address_next<= 106 ;
        2013 : Address_next<= 107 ;
        2014 : Address_next<= 214 ;
        2015 : Address_next<= 428 ;
        2017 : Address_next<= 429 ;
        2018 : Address_next<= 214 ;
        2020 : Address_next<= 215 ;
        2021 : Address_next<= 430 ;
        2023 : Address_next<= 431 ;
        2024 : Address_next<= 215 ;
        2025 : Address_next<= 107 ;
        2026 : Address_next<= 53 ;
        2027 : Address_next<= 26 ;
        2030 : Address_next<= 27 ;
        2031 : Address_next<= 54 ;
        2032 : Address_next<= 108 ;
        2033 : Address_next<= 216 ;
        2034 : Address_next<= 432 ;
        2036 : Address_next<= 433 ;
        2037 : Address_next<= 216 ;
        2039 : Address_next<= 217 ;
        2040 : Address_next<= 434 ;
        2042 : Address_next<= 435 ;
        2043 : Address_next<= 217 ;
        2044 : Address_next<= 108 ;
        2046 : Address_next<= 109 ;
        2047 : Address_next<= 218 ;
        2048 : Address_next<= 436 ;
        2050 : Address_next<= 437 ;
        2051 : Address_next<= 218 ;
        2053 : Address_next<= 219 ;
        2054 : Address_next<= 438 ;
        2056 : Address_next<= 439 ;
        2057 : Address_next<= 219 ;
        2058 : Address_next<= 109 ;
        2059 : Address_next<= 54 ;
        2061 : Address_next<= 55 ;
        2062 : Address_next<= 110 ;
        2063 : Address_next<= 220 ;
        2064 : Address_next<= 440 ;
        2066 : Address_next<= 441 ;
        2067 : Address_next<= 220 ;
        2069 : Address_next<= 221 ;
        2070 : Address_next<= 442 ;
        2072 : Address_next<= 443 ;
        2073 : Address_next<= 221 ;
        2074 : Address_next<= 110 ;
        2076 : Address_next<= 111 ;
        2077 : Address_next<= 222 ;
        2078 : Address_next<= 444 ;
        2080 : Address_next<= 445 ;
        2081 : Address_next<= 222 ;
        2083 : Address_next<= 223 ;
        2084 : Address_next<= 446 ;
        2086 : Address_next<= 447 ;
        2087 : Address_next<= 223 ;
        2088 : Address_next<= 111 ;
        2089 : Address_next<= 55 ;
        2090 : Address_next<= 27 ;
        2091 : Address_next<= 13 ;
        2092 : Address_next<= 13 ;
        2093 : Address_next<= 6 ;
        2094 : Address_next<= 6 ;
        2095 : Address_next<= 6 ;
        2096 : Address_next<= 6 ;
        2105 : Address_next<= 7 ;
        2106 : Address_next<= 7 ;
        2107 : Address_next<= 7 ;
        2108 : Address_next<= 7 ;
        2109 : Address_next<= 14 ;
        2110 : Address_next<= 14 ;
        2111 : Address_next<= 28 ;
        2112 : Address_next<= 56 ;
        2113 : Address_next<= 112 ;
        2114 : Address_next<= 224 ;
        2115 : Address_next<= 448 ;
        2117 : Address_next<= 449 ;
        2118 : Address_next<= 224 ;
        2120 : Address_next<= 225 ;
        2121 : Address_next<= 450 ;
        2123 : Address_next<= 451 ;
        2124 : Address_next<= 225 ;
        2125 : Address_next<= 112 ;
        2127 : Address_next<= 113 ;
        2128 : Address_next<= 226 ;
        2129 : Address_next<= 452 ;
        2131 : Address_next<= 453 ;
        2132 : Address_next<= 226 ;
        2134 : Address_next<= 227 ;
        2135 : Address_next<= 454 ;
        2137 : Address_next<= 455 ;
        2138 : Address_next<= 227 ;
        2139 : Address_next<= 113 ;
        2140 : Address_next<= 56 ;
        2142 : Address_next<= 57 ;
        2143 : Address_next<= 114 ;
        2144 : Address_next<= 228 ;
        2145 : Address_next<= 456 ;
        2147 : Address_next<= 457 ;
        2148 : Address_next<= 228 ;
        2150 : Address_next<= 229 ;
        2151 : Address_next<= 458 ;
        2153 : Address_next<= 459 ;
        2154 : Address_next<= 229 ;
        2155 : Address_next<= 114 ;
        2157 : Address_next<= 115 ;
        2158 : Address_next<= 230 ;
        2159 : Address_next<= 460 ;
        2161 : Address_next<= 461 ;
        2162 : Address_next<= 230 ;
        2164 : Address_next<= 231 ;
        2165 : Address_next<= 462 ;
        2167 : Address_next<= 463 ;
        2168 : Address_next<= 231 ;
        2169 : Address_next<= 115 ;
        2170 : Address_next<= 57 ;
        2171 : Address_next<= 28 ;
        2174 : Address_next<= 29 ;
        2175 : Address_next<= 58 ;
        2176 : Address_next<= 116 ;
        2177 : Address_next<= 232 ;
        2178 : Address_next<= 464 ;
        2180 : Address_next<= 465 ;
        2181 : Address_next<= 232 ;
        2183 : Address_next<= 233 ;
        2184 : Address_next<= 466 ;
        2186 : Address_next<= 467 ;
        2187 : Address_next<= 233 ;
        2188 : Address_next<= 116 ;
        2190 : Address_next<= 117 ;
        2191 : Address_next<= 234 ;
        2192 : Address_next<= 468 ;
        2194 : Address_next<= 469 ;
        2195 : Address_next<= 234 ;
        2197 : Address_next<= 235 ;
        2198 : Address_next<= 470 ;
        2200 : Address_next<= 471 ;
        2201 : Address_next<= 235 ;
        2202 : Address_next<= 117 ;
        2203 : Address_next<= 58 ;
        2205 : Address_next<= 59 ;
        2206 : Address_next<= 118 ;
        2207 : Address_next<= 236 ;
        2208 : Address_next<= 472 ;
        2210 : Address_next<= 473 ;
        2211 : Address_next<= 236 ;
        2213 : Address_next<= 237 ;
        2214 : Address_next<= 474 ;
        2216 : Address_next<= 475 ;
        2217 : Address_next<= 237 ;
        2218 : Address_next<= 118 ;
        2220 : Address_next<= 119 ;
        2221 : Address_next<= 238 ;
        2222 : Address_next<= 476 ;
        2224 : Address_next<= 477 ;
        2225 : Address_next<= 238 ;
        2227 : Address_next<= 239 ;
        2228 : Address_next<= 478 ;
        2230 : Address_next<= 479 ;
        2231 : Address_next<= 239 ;
        2232 : Address_next<= 119 ;
        2233 : Address_next<= 59 ;
        2234 : Address_next<= 29 ;
        2235 : Address_next<= 14 ;
        2236 : Address_next<= 14 ;
        2241 : Address_next<= 15 ;
        2242 : Address_next<= 15 ;
        2243 : Address_next<= 30 ;
        2244 : Address_next<= 60 ;
        2245 : Address_next<= 120 ;
        2246 : Address_next<= 240 ;
        2247 : Address_next<= 480 ;
        2249 : Address_next<= 481 ;
        2250 : Address_next<= 240 ;
        2252 : Address_next<= 241 ;
        2253 : Address_next<= 482 ;
        2255 : Address_next<= 483 ;
        2256 : Address_next<= 241 ;
        2257 : Address_next<= 120 ;
        2259 : Address_next<= 121 ;
        2260 : Address_next<= 242 ;
        2261 : Address_next<= 484 ;
        2263 : Address_next<= 485 ;
        2264 : Address_next<= 242 ;
        2266 : Address_next<= 243 ;
        2267 : Address_next<= 486 ;
        2269 : Address_next<= 487 ;
        2270 : Address_next<= 243 ;
        2271 : Address_next<= 121 ;
        2272 : Address_next<= 60 ;
        2274 : Address_next<= 61 ;
        2275 : Address_next<= 122 ;
        2276 : Address_next<= 244 ;
        2277 : Address_next<= 488 ;
        2279 : Address_next<= 489 ;
        2280 : Address_next<= 244 ;
        2282 : Address_next<= 245 ;
        2283 : Address_next<= 490 ;
        2285 : Address_next<= 491 ;
        2286 : Address_next<= 245 ;
        2287 : Address_next<= 122 ;
        2289 : Address_next<= 123 ;
        2290 : Address_next<= 246 ;
        2291 : Address_next<= 492 ;
        2293 : Address_next<= 493 ;
        2294 : Address_next<= 246 ;
        2296 : Address_next<= 247 ;
        2297 : Address_next<= 494 ;
        2299 : Address_next<= 495 ;
        2300 : Address_next<= 247 ;
        2301 : Address_next<= 123 ;
        2302 : Address_next<= 61 ;
        2303 : Address_next<= 30 ;
        2306 : Address_next<= 31 ;
        2307 : Address_next<= 62 ;
        2308 : Address_next<= 124 ;
        2309 : Address_next<= 248 ;
        2310 : Address_next<= 496 ;
        2312 : Address_next<= 497 ;
        2313 : Address_next<= 248 ;
        2315 : Address_next<= 249 ;
        2316 : Address_next<= 498 ;
        2318 : Address_next<= 499 ;
        2319 : Address_next<= 249 ;
        2320 : Address_next<= 124 ;
        2322 : Address_next<= 125 ;
        2323 : Address_next<= 250 ;
        2324 : Address_next<= 500 ;
        2326 : Address_next<= 501 ;
        2327 : Address_next<= 250 ;
        2329 : Address_next<= 251 ;
        2330 : Address_next<= 502 ;
        2332 : Address_next<= 503 ;
        2333 : Address_next<= 251 ;
        2334 : Address_next<= 125 ;
        2335 : Address_next<= 62 ;
        2337 : Address_next<= 63 ;
        2338 : Address_next<= 126 ;
        2339 : Address_next<= 252 ;
        2340 : Address_next<= 504 ;
        2342 : Address_next<= 505 ;
        2343 : Address_next<= 252 ;
        2345 : Address_next<= 253 ;
        2346 : Address_next<= 506 ;
        2348 : Address_next<= 507 ;
        2349 : Address_next<= 253 ;
        2350 : Address_next<= 126 ;
        2352 : Address_next<= 127 ;
        2353 : Address_next<= 254 ;
        2354 : Address_next<= 508 ;
        2356 : Address_next<= 509 ;
        2357 : Address_next<= 254 ;
        2359 : Address_next<= 255 ;
        2360 : Address_next<= 510 ;
        2362 : Address_next<= 511 ;
        2363 : Address_next<= 255 ;
        2364 : Address_next<= 127 ;
        2365 : Address_next<= 63 ;
        2366 : Address_next<= 31 ;
        2367 : Address_next<= 15 ;
        2368 : Address_next<= 15 ;
        2369 : Address_next<= 7 ;
        2370 : Address_next<= 7 ;
        2371 : Address_next<= 7 ;
        2372 : Address_next<= 7 ;
        2373 : Address_next<= 3 ;
        2374 : Address_next<= 3 ;
        2375 : Address_next<= 3 ;
        2376 : Address_next<= 3 ;
        2377 : Address_next<= 3 ;
        2378 : Address_next<= 3 ;
        2379 : Address_next<= 3 ;
        2380 : Address_next<= 3 ;
        2381 : Address_next<= 1 ;
        2382 : Address_next<= 1 ;
        2383 : Address_next<= 1 ;
        2384 : Address_next<= 1 ;
        2385 : Address_next<= 1 ;
        2386 : Address_next<= 1 ;
        2387 : Address_next<= 1 ;
        2388 : Address_next<= 1 ;
        2389 : Address_next<= 1 ;
        2390 : Address_next<= 1 ;
        2391 : Address_next<= 1 ;
        2392 : Address_next<= 1 ;
        2393 : Address_next<= 1 ;
        2394 : Address_next<= 1 ;
        2395 : Address_next<= 1 ;
        2396 : Address_next<= 1 ;
        default : Address_next <= 0;
       endcase

      end
      else begin
           L_Nv_next                     <=1024;
           L_opcode_next <= TYPE1;
           L_part_count_next <= 0;
           Address_next <= 0;
      end
end
end
endmodule


